// This is the unpowered netlist.
module cawb (ca_dbus_ack,
    ca_dbus_com,
    ca_dbus_valid,
    ca_match_ack,
    ca_match_valid,
    ca_time_ack,
    ca_time_valid,
    cubev_ca_clk0,
    cubev_ca_clk1,
    cubev_ca_csb0,
    cubev_ca_csb1,
    cubev_ca_web0,
    cubev_phi_clk0,
    cubev_phi_csb0,
    cubev_phi_web0,
    cubev_pli_clk0,
    cubev_pli_csb0,
    cubev_pli_web0,
    rstn_reg,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    ca_command,
    ca_dbus_data,
    ca_dbus_tid,
    ca_time_data,
    cubev_ca_addr0,
    cubev_ca_addr1,
    cubev_ca_din0,
    cubev_ca_dout0,
    cubev_ca_dout1,
    cubev_ca_wmask0,
    cubev_phi_addr0,
    cubev_phi_din0,
    cubev_phi_dout0,
    cubev_phi_wmask0,
    cubev_pli_addr0,
    cubev_pli_din0,
    cubev_pli_dout0,
    cubev_pli_wmask0,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 output ca_dbus_ack;
 input ca_dbus_com;
 input ca_dbus_valid;
 input ca_match_ack;
 output ca_match_valid;
 input ca_time_ack;
 output ca_time_valid;
 output cubev_ca_clk0;
 output cubev_ca_clk1;
 output cubev_ca_csb0;
 output cubev_ca_csb1;
 output cubev_ca_web0;
 output cubev_phi_clk0;
 output cubev_phi_csb0;
 output cubev_phi_web0;
 output cubev_pli_clk0;
 output cubev_pli_csb0;
 output cubev_pli_web0;
 output rstn_reg;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [31:0] ca_command;
 input [31:0] ca_dbus_data;
 input [2:0] ca_dbus_tid;
 output [22:0] ca_time_data;
 output [7:0] cubev_ca_addr0;
 output [7:0] cubev_ca_addr1;
 output [31:0] cubev_ca_din0;
 input [31:0] cubev_ca_dout0;
 input [31:0] cubev_ca_dout1;
 output [3:0] cubev_ca_wmask0;
 output [7:0] cubev_phi_addr0;
 output [31:0] cubev_phi_din0;
 input [31:0] cubev_phi_dout0;
 output [3:0] cubev_phi_wmask0;
 output [7:0] cubev_pli_addr0;
 output [31:0] cubev_pli_din0;
 input [31:0] cubev_pli_dout0;
 output [3:0] cubev_pli_wmask0;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire net755;
 wire _0074_;
 wire net756;
 wire _0076_;
 wire net757;
 wire _0078_;
 wire net758;
 wire _0080_;
 wire net759;
 wire _0082_;
 wire net760;
 wire _0084_;
 wire net761;
 wire _0086_;
 wire net762;
 wire _0088_;
 wire net763;
 wire _0090_;
 wire net764;
 wire _0092_;
 wire net765;
 wire _0094_;
 wire net766;
 wire _0096_;
 wire net767;
 wire _0098_;
 wire net768;
 wire _0100_;
 wire net769;
 wire _0102_;
 wire net770;
 wire _0104_;
 wire net771;
 wire _0106_;
 wire net772;
 wire _0108_;
 wire net773;
 wire _0110_;
 wire net774;
 wire _0112_;
 wire net775;
 wire _0114_;
 wire net776;
 wire _0116_;
 wire net777;
 wire _0118_;
 wire net778;
 wire _0120_;
 wire net779;
 wire _0122_;
 wire net780;
 wire _0124_;
 wire net781;
 wire _0126_;
 wire net782;
 wire _0128_;
 wire net783;
 wire _0130_;
 wire net784;
 wire _0132_;
 wire net785;
 wire _0134_;
 wire net786;
 wire _0136_;
 wire net787;
 wire _0138_;
 wire net788;
 wire _0140_;
 wire net789;
 wire _0142_;
 wire net790;
 wire _0144_;
 wire net791;
 wire _0146_;
 wire net792;
 wire _0148_;
 wire net793;
 wire _0150_;
 wire net794;
 wire _0152_;
 wire net795;
 wire _0154_;
 wire net796;
 wire _0156_;
 wire net797;
 wire _0158_;
 wire net798;
 wire _0160_;
 wire net799;
 wire _0162_;
 wire net800;
 wire _0164_;
 wire net801;
 wire _0166_;
 wire net802;
 wire _0168_;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire _0202_;
 wire net836;
 wire _0204_;
 wire net837;
 wire _0206_;
 wire net838;
 wire _0208_;
 wire net839;
 wire _0210_;
 wire net840;
 wire _0212_;
 wire net841;
 wire _0214_;
 wire net842;
 wire _0216_;
 wire net843;
 wire _0218_;
 wire net844;
 wire _0220_;
 wire net845;
 wire _0222_;
 wire net846;
 wire _0224_;
 wire net847;
 wire _0226_;
 wire net848;
 wire _0228_;
 wire net849;
 wire _0230_;
 wire net850;
 wire _0232_;
 wire net851;
 wire _0234_;
 wire net852;
 wire _0236_;
 wire net853;
 wire _0238_;
 wire net854;
 wire _0240_;
 wire net855;
 wire _0242_;
 wire net856;
 wire _0244_;
 wire net857;
 wire _0246_;
 wire net858;
 wire _0248_;
 wire net859;
 wire _0250_;
 wire net860;
 wire _0252_;
 wire net861;
 wire _0254_;
 wire net862;
 wire _0256_;
 wire net863;
 wire _0258_;
 wire net864;
 wire _0260_;
 wire net865;
 wire _0262_;
 wire net866;
 wire _0264_;
 wire net867;
 wire _0266_;
 wire net868;
 wire _0268_;
 wire net869;
 wire _0270_;
 wire net870;
 wire _0272_;
 wire net871;
 wire _0274_;
 wire net872;
 wire _0276_;
 wire net873;
 wire _0278_;
 wire clknet_leaf_1_wb_clk_i;
 wire _0280_;
 wire net695;
 wire _0282_;
 wire net696;
 wire _0284_;
 wire net697;
 wire _0286_;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire net634;
 wire net635;
 wire net636;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net637;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net638;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire \i_ca.ca_compare_check ;
 wire \i_ca.ca_dbus_valid_meta ;
 wire \i_ca.ca_end_of_wr_list ;
 wire \i_ca.ca_insert_equal_high ;
 wire \i_ca.ca_insert_lesser_high ;
 wire \i_ca.ca_insert_lesser_low ;
 wire \i_ca.ca_insert_time[0] ;
 wire \i_ca.ca_insert_time[10] ;
 wire \i_ca.ca_insert_time[11] ;
 wire \i_ca.ca_insert_time[12] ;
 wire \i_ca.ca_insert_time[13] ;
 wire \i_ca.ca_insert_time[14] ;
 wire \i_ca.ca_insert_time[15] ;
 wire \i_ca.ca_insert_time[16] ;
 wire \i_ca.ca_insert_time[17] ;
 wire \i_ca.ca_insert_time[18] ;
 wire \i_ca.ca_insert_time[19] ;
 wire \i_ca.ca_insert_time[1] ;
 wire \i_ca.ca_insert_time[20] ;
 wire \i_ca.ca_insert_time[21] ;
 wire \i_ca.ca_insert_time[22] ;
 wire \i_ca.ca_insert_time[2] ;
 wire \i_ca.ca_insert_time[3] ;
 wire \i_ca.ca_insert_time[4] ;
 wire \i_ca.ca_insert_time[5] ;
 wire \i_ca.ca_insert_time[6] ;
 wire \i_ca.ca_insert_time[7] ;
 wire \i_ca.ca_insert_time[8] ;
 wire \i_ca.ca_insert_time[9] ;
 wire \i_ca.ca_match_ack_meta ;
 wire \i_ca.ca_match_block_ack ;
 wire \i_ca.ca_match_check ;
 wire \i_ca.ca_match_hs_state[0] ;
 wire \i_ca.ca_match_hs_state[1] ;
 wire \i_ca.ca_match_hs_state[2] ;
 wire \i_ca.ca_match_req ;
 wire \i_ca.ca_rd_add[0] ;
 wire \i_ca.ca_rd_add[1] ;
 wire \i_ca.ca_rd_add[2] ;
 wire \i_ca.ca_rd_add[3] ;
 wire \i_ca.ca_rd_add[4] ;
 wire \i_ca.ca_rd_add[5] ;
 wire \i_ca.ca_rd_add[6] ;
 wire \i_ca.ca_rd_add[7] ;
 wire \i_ca.ca_rd_doutb[0] ;
 wire \i_ca.ca_rd_doutb[10] ;
 wire \i_ca.ca_rd_doutb[11] ;
 wire \i_ca.ca_rd_doutb[12] ;
 wire \i_ca.ca_rd_doutb[13] ;
 wire \i_ca.ca_rd_doutb[14] ;
 wire \i_ca.ca_rd_doutb[15] ;
 wire \i_ca.ca_rd_doutb[16] ;
 wire \i_ca.ca_rd_doutb[17] ;
 wire \i_ca.ca_rd_doutb[18] ;
 wire \i_ca.ca_rd_doutb[19] ;
 wire \i_ca.ca_rd_doutb[1] ;
 wire \i_ca.ca_rd_doutb[20] ;
 wire \i_ca.ca_rd_doutb[21] ;
 wire \i_ca.ca_rd_doutb[22] ;
 wire \i_ca.ca_rd_doutb[23] ;
 wire \i_ca.ca_rd_doutb[24] ;
 wire \i_ca.ca_rd_doutb[25] ;
 wire \i_ca.ca_rd_doutb[26] ;
 wire \i_ca.ca_rd_doutb[27] ;
 wire \i_ca.ca_rd_doutb[28] ;
 wire \i_ca.ca_rd_doutb[29] ;
 wire \i_ca.ca_rd_doutb[2] ;
 wire \i_ca.ca_rd_doutb[30] ;
 wire \i_ca.ca_rd_doutb[32] ;
 wire \i_ca.ca_rd_doutb[3] ;
 wire \i_ca.ca_rd_doutb[4] ;
 wire \i_ca.ca_rd_doutb[5] ;
 wire \i_ca.ca_rd_doutb[6] ;
 wire \i_ca.ca_rd_doutb[7] ;
 wire \i_ca.ca_rd_doutb[8] ;
 wire \i_ca.ca_rd_doutb[9] ;
 wire \i_ca.ca_rd_doutb_31_23 ;
 wire \i_ca.ca_rd_doutb_32 ;
 wire \i_ca.ca_rd_fsm_state[0] ;
 wire \i_ca.ca_rd_fsm_state[1] ;
 wire \i_ca.ca_rd_fsm_state[2] ;
 wire \i_ca.ca_rd_fsm_state[3] ;
 wire \i_ca.ca_rd_fsm_state[4] ;
 wire \i_ca.ca_rd_fsm_state[5] ;
 wire \i_ca.ca_rd_fsm_state[6] ;
 wire \i_ca.ca_rd_fsm_state[7] ;
 wire \i_ca.ca_rd_fsm_state[8] ;
 wire \i_ca.ca_ready ;
 wire \i_ca.ca_time_const[0] ;
 wire \i_ca.ca_time_const[10] ;
 wire \i_ca.ca_time_const[11] ;
 wire \i_ca.ca_time_const[12] ;
 wire \i_ca.ca_time_const[13] ;
 wire \i_ca.ca_time_const[14] ;
 wire \i_ca.ca_time_const[15] ;
 wire \i_ca.ca_time_const[16] ;
 wire \i_ca.ca_time_const[17] ;
 wire \i_ca.ca_time_const[18] ;
 wire \i_ca.ca_time_const[19] ;
 wire \i_ca.ca_time_const[1] ;
 wire \i_ca.ca_time_const[20] ;
 wire \i_ca.ca_time_const[21] ;
 wire \i_ca.ca_time_const[22] ;
 wire \i_ca.ca_time_const[2] ;
 wire \i_ca.ca_time_const[3] ;
 wire \i_ca.ca_time_const[4] ;
 wire \i_ca.ca_time_const[5] ;
 wire \i_ca.ca_time_const[6] ;
 wire \i_ca.ca_time_const[7] ;
 wire \i_ca.ca_time_const[8] ;
 wire \i_ca.ca_time_const[9] ;
 wire \i_ca.ca_time_diff[12] ;
 wire \i_ca.ca_time_diff[13] ;
 wire \i_ca.ca_time_diff[14] ;
 wire \i_ca.ca_time_diff[15] ;
 wire \i_ca.ca_time_diff[16] ;
 wire \i_ca.ca_time_diff[17] ;
 wire \i_ca.ca_time_diff[18] ;
 wire \i_ca.ca_time_diff[19] ;
 wire \i_ca.ca_time_diff[20] ;
 wire \i_ca.ca_time_diff[21] ;
 wire \i_ca.ca_time_diff[22] ;
 wire \i_ca.ca_update_rd_add ;
 wire \i_ca.ca_wr_add[0] ;
 wire \i_ca.ca_wr_add[1] ;
 wire \i_ca.ca_wr_add[2] ;
 wire \i_ca.ca_wr_add[3] ;
 wire \i_ca.ca_wr_add[4] ;
 wire \i_ca.ca_wr_add[5] ;
 wire \i_ca.ca_wr_add[6] ;
 wire \i_ca.ca_wr_add[7] ;
 wire \i_ca.ca_wr_add[8] ;
 wire \i_ca.ca_wr_add_fill[1] ;
 wire \i_ca.ca_wr_add_fill[2] ;
 wire \i_ca.ca_wr_add_fill[3] ;
 wire \i_ca.ca_wr_add_fill[4] ;
 wire \i_ca.ca_wr_add_fill[5] ;
 wire \i_ca.ca_wr_add_fill[6] ;
 wire \i_ca.ca_wr_add_fill[7] ;
 wire \i_ca.ca_wr_add_fill[8] ;
 wire \i_ca.ca_wr_add_ptr[0] ;
 wire \i_ca.ca_wr_add_ptr[1] ;
 wire \i_ca.ca_wr_add_ptr[2] ;
 wire \i_ca.ca_wr_add_ptr[3] ;
 wire \i_ca.ca_wr_add_ptr[4] ;
 wire \i_ca.ca_wr_add_ptr[5] ;
 wire \i_ca.ca_wr_add_ptr[6] ;
 wire \i_ca.ca_wr_add_ptr[7] ;
 wire \i_ca.ca_wr_add_ptr[8] ;
 wire \i_ca.ca_wr_add_start[0] ;
 wire \i_ca.ca_wr_add_start[1] ;
 wire \i_ca.ca_wr_add_start[2] ;
 wire \i_ca.ca_wr_add_start[3] ;
 wire \i_ca.ca_wr_add_start[4] ;
 wire \i_ca.ca_wr_add_start[5] ;
 wire \i_ca.ca_wr_add_start[6] ;
 wire \i_ca.ca_wr_add_start[7] ;
 wire \i_ca.ca_wr_add_start[8] ;
 wire \i_ca.ca_wr_add_start_marker ;
 wire \i_ca.ca_wr_com_const ;
 wire \i_ca.ca_wr_dina[0] ;
 wire \i_ca.ca_wr_dina[10] ;
 wire \i_ca.ca_wr_dina[11] ;
 wire \i_ca.ca_wr_dina[12] ;
 wire \i_ca.ca_wr_dina[13] ;
 wire \i_ca.ca_wr_dina[14] ;
 wire \i_ca.ca_wr_dina[15] ;
 wire \i_ca.ca_wr_dina[16] ;
 wire \i_ca.ca_wr_dina[17] ;
 wire \i_ca.ca_wr_dina[18] ;
 wire \i_ca.ca_wr_dina[19] ;
 wire \i_ca.ca_wr_dina[1] ;
 wire \i_ca.ca_wr_dina[20] ;
 wire \i_ca.ca_wr_dina[21] ;
 wire \i_ca.ca_wr_dina[22] ;
 wire \i_ca.ca_wr_dina[23] ;
 wire \i_ca.ca_wr_dina[24] ;
 wire \i_ca.ca_wr_dina[25] ;
 wire \i_ca.ca_wr_dina[26] ;
 wire \i_ca.ca_wr_dina[27] ;
 wire \i_ca.ca_wr_dina[28] ;
 wire \i_ca.ca_wr_dina[29] ;
 wire \i_ca.ca_wr_dina[2] ;
 wire \i_ca.ca_wr_dina[30] ;
 wire \i_ca.ca_wr_dina[31] ;
 wire \i_ca.ca_wr_dina[32] ;
 wire \i_ca.ca_wr_dina[3] ;
 wire \i_ca.ca_wr_dina[4] ;
 wire \i_ca.ca_wr_dina[5] ;
 wire \i_ca.ca_wr_dina[6] ;
 wire \i_ca.ca_wr_dina[7] ;
 wire \i_ca.ca_wr_dina[8] ;
 wire \i_ca.ca_wr_dina[9] ;
 wire \i_ca.ca_wr_douta[0] ;
 wire \i_ca.ca_wr_douta[10] ;
 wire \i_ca.ca_wr_douta[11] ;
 wire \i_ca.ca_wr_douta[12] ;
 wire \i_ca.ca_wr_douta[13] ;
 wire \i_ca.ca_wr_douta[14] ;
 wire \i_ca.ca_wr_douta[15] ;
 wire \i_ca.ca_wr_douta[16] ;
 wire \i_ca.ca_wr_douta[17] ;
 wire \i_ca.ca_wr_douta[18] ;
 wire \i_ca.ca_wr_douta[19] ;
 wire \i_ca.ca_wr_douta[1] ;
 wire \i_ca.ca_wr_douta[20] ;
 wire \i_ca.ca_wr_douta[21] ;
 wire \i_ca.ca_wr_douta[22] ;
 wire \i_ca.ca_wr_douta[23] ;
 wire \i_ca.ca_wr_douta[24] ;
 wire \i_ca.ca_wr_douta[25] ;
 wire \i_ca.ca_wr_douta[26] ;
 wire \i_ca.ca_wr_douta[27] ;
 wire \i_ca.ca_wr_douta[28] ;
 wire \i_ca.ca_wr_douta[29] ;
 wire \i_ca.ca_wr_douta[2] ;
 wire \i_ca.ca_wr_douta[30] ;
 wire \i_ca.ca_wr_douta[32] ;
 wire \i_ca.ca_wr_douta[3] ;
 wire \i_ca.ca_wr_douta[4] ;
 wire \i_ca.ca_wr_douta[5] ;
 wire \i_ca.ca_wr_douta[6] ;
 wire \i_ca.ca_wr_douta[7] ;
 wire \i_ca.ca_wr_douta[8] ;
 wire \i_ca.ca_wr_douta[9] ;
 wire \i_ca.ca_wr_et_const ;
 wire \i_ca.ca_wr_fsm_state[0] ;
 wire \i_ca.ca_wr_fsm_state[10] ;
 wire \i_ca.ca_wr_fsm_state[11] ;
 wire \i_ca.ca_wr_fsm_state[12] ;
 wire \i_ca.ca_wr_fsm_state[13] ;
 wire \i_ca.ca_wr_fsm_state[14] ;
 wire \i_ca.ca_wr_fsm_state[15] ;
 wire \i_ca.ca_wr_fsm_state[16] ;
 wire \i_ca.ca_wr_fsm_state[17] ;
 wire \i_ca.ca_wr_fsm_state[1] ;
 wire \i_ca.ca_wr_fsm_state[2] ;
 wire \i_ca.ca_wr_fsm_state[3] ;
 wire \i_ca.ca_wr_fsm_state[4] ;
 wire \i_ca.ca_wr_fsm_state[5] ;
 wire \i_ca.ca_wr_fsm_state[6] ;
 wire \i_ca.ca_wr_fsm_state[7] ;
 wire \i_ca.ca_wr_fsm_state[8] ;
 wire \i_ca.ca_wr_fsm_state[9] ;
 wire \i_ca.ca_wr_sync_update ;
 wire \i_ca.ca_wr_sync_update_done ;
 wire \i_ca.ca_wr_wea ;
 wire \i_ca.cubev_ca_wea ;
 wire \i_ca.hs_ready_meta ;
 wire \i_ca.hs_state_write_const[0] ;
 wire \i_ca.hs_state_write_const[1] ;
 wire \i_ca.hs_state_write_const[2] ;
 wire \i_ca.hs_state_write_const[3] ;
 wire \i_ca.hs_write_dbus_wr_data_const[0] ;
 wire \i_ca.hs_write_dbus_wr_data_const[10] ;
 wire \i_ca.hs_write_dbus_wr_data_const[11] ;
 wire \i_ca.hs_write_dbus_wr_data_const[12] ;
 wire \i_ca.hs_write_dbus_wr_data_const[13] ;
 wire \i_ca.hs_write_dbus_wr_data_const[14] ;
 wire \i_ca.hs_write_dbus_wr_data_const[15] ;
 wire \i_ca.hs_write_dbus_wr_data_const[16] ;
 wire \i_ca.hs_write_dbus_wr_data_const[17] ;
 wire \i_ca.hs_write_dbus_wr_data_const[18] ;
 wire \i_ca.hs_write_dbus_wr_data_const[19] ;
 wire \i_ca.hs_write_dbus_wr_data_const[1] ;
 wire \i_ca.hs_write_dbus_wr_data_const[20] ;
 wire \i_ca.hs_write_dbus_wr_data_const[21] ;
 wire \i_ca.hs_write_dbus_wr_data_const[22] ;
 wire \i_ca.hs_write_dbus_wr_data_const[23] ;
 wire \i_ca.hs_write_dbus_wr_data_const[24] ;
 wire \i_ca.hs_write_dbus_wr_data_const[25] ;
 wire \i_ca.hs_write_dbus_wr_data_const[26] ;
 wire \i_ca.hs_write_dbus_wr_data_const[27] ;
 wire \i_ca.hs_write_dbus_wr_data_const[28] ;
 wire \i_ca.hs_write_dbus_wr_data_const[29] ;
 wire \i_ca.hs_write_dbus_wr_data_const[2] ;
 wire \i_ca.hs_write_dbus_wr_data_const[30] ;
 wire \i_ca.hs_write_dbus_wr_data_const[31] ;
 wire \i_ca.hs_write_dbus_wr_data_const[3] ;
 wire \i_ca.hs_write_dbus_wr_data_const[4] ;
 wire \i_ca.hs_write_dbus_wr_data_const[5] ;
 wire \i_ca.hs_write_dbus_wr_data_const[6] ;
 wire \i_ca.hs_write_dbus_wr_data_const[7] ;
 wire \i_ca.hs_write_dbus_wr_data_const[8] ;
 wire \i_ca.hs_write_dbus_wr_data_const[9] ;
 wire \i_ca.hs_write_tid_wr0_const[0] ;
 wire \i_ca.hs_write_tid_wr0_const[1] ;
 wire \i_ca.hs_write_tid_wr0_const[2] ;
 wire net639;
 wire net640;
 wire net641;
 wire net673;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire prog_h_addr0;
 wire prog_wea;
 wire net674;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0_0_wb_clk_i;
 wire clknet_1_0_1_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_1_1_1_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_2_1_wb_clk_i;
 wire clknet_opt_2_2_wb_clk_i;
 wire clknet_opt_2_3_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_3_1_wb_clk_i;
 wire clknet_opt_3_2_wb_clk_i;
 wire clknet_opt_4_0_wb_clk_i;
 wire clknet_opt_4_1_wb_clk_i;
 wire clknet_opt_5_0_wb_clk_i;
 wire clknet_0__0983_;
 wire clknet_1_0__leaf__0983_;
 wire clknet_1_1__leaf__0983_;
 wire clknet_0__1029_;
 wire clknet_1_0__leaf__1029_;
 wire clknet_1_1__leaf__1029_;
 wire clknet_0__1028_;
 wire clknet_1_0__leaf__1028_;
 wire clknet_1_1__leaf__1028_;
 wire clknet_0__1027_;
 wire clknet_1_0__leaf__1027_;
 wire clknet_1_1__leaf__1027_;
 wire clknet_0__1026_;
 wire clknet_1_0__leaf__1026_;
 wire clknet_1_1__leaf__1026_;
 wire clknet_0__1025_;
 wire clknet_1_0__leaf__1025_;
 wire clknet_1_1__leaf__1025_;
 wire clknet_0__1024_;
 wire clknet_1_0__leaf__1024_;
 wire clknet_1_1__leaf__1024_;
 wire clknet_0__0987_;
 wire clknet_1_0_0__0987_;
 wire clknet_1_1_0__0987_;
 wire clknet_0__1023_;
 wire clknet_1_0__leaf__1023_;
 wire clknet_1_1__leaf__1023_;
 wire clknet_0__1022_;
 wire clknet_1_0__leaf__1022_;
 wire clknet_1_1__leaf__1022_;
 wire clknet_0__1021_;
 wire clknet_1_0__leaf__1021_;
 wire clknet_1_1__leaf__1021_;
 wire clknet_0__0994_;
 wire clknet_1_0__leaf__0994_;
 wire clknet_1_1__leaf__0994_;
 wire clknet_0__0993_;
 wire clknet_1_0__leaf__0993_;
 wire clknet_1_1__leaf__0993_;
 wire clknet_0__0992_;
 wire clknet_1_0__leaf__0992_;
 wire clknet_1_1__leaf__0992_;
 wire clknet_0__0991_;
 wire clknet_1_0__leaf__0991_;
 wire clknet_1_1__leaf__0991_;
 wire clknet_0__0990_;
 wire clknet_1_0__leaf__0990_;
 wire clknet_1_1__leaf__0990_;
 wire clknet_0__0989_;
 wire clknet_1_0__leaf__0989_;
 wire clknet_1_1__leaf__0989_;
 wire clknet_0__0988_;
 wire clknet_1_0__leaf__0988_;
 wire clknet_1_1__leaf__0988_;
 wire clknet_0__0984_;
 wire clknet_1_0__leaf__0984_;
 wire clknet_1_1__leaf__0984_;
 wire clknet_0__0986_;
 wire clknet_1_0__leaf__0986_;
 wire clknet_1_1__leaf__0986_;
 wire clknet_0__0985_;
 wire clknet_1_0__leaf__0985_;
 wire clknet_1_1__leaf__0985_;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;

 sky130_fd_sc_hd__buf_12 _1439_ (.A(net211),
    .X(_0589_));
 sky130_fd_sc_hd__buf_6 _1440_ (.A(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__inv_2 _1441_ (.A(_0590_),
    .Y(_0286_));
 sky130_fd_sc_hd__buf_4 _1442_ (.A(net205),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _1443_ (.A0(net265),
    .A1(net192),
    .S(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__inv_2 _1444_ (.A(net205),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(net273),
    .B(net240),
    .Y(_0594_));
 sky130_fd_sc_hd__or4_1 _1446_ (.A(net216),
    .B(net217),
    .C(net220),
    .D(net223),
    .X(_0595_));
 sky130_fd_sc_hd__or4b_1 _1447_ (.A(net224),
    .B(net227),
    .C(net231),
    .D_N(net228),
    .X(_0596_));
 sky130_fd_sc_hd__or4_1 _1448_ (.A(net215),
    .B(net218),
    .C(net221),
    .D(net222),
    .X(_0597_));
 sky130_fd_sc_hd__or4b_1 _1449_ (.A(net225),
    .B(net226),
    .C(net232),
    .D_N(net229),
    .X(_0598_));
 sky130_fd_sc_hd__or4_2 _1450_ (.A(_0595_),
    .B(_0596_),
    .C(_0597_),
    .D(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or4b_2 _1451_ (.A(net206),
    .B(_0594_),
    .C(_0599_),
    .D_N(net274),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_4 _1452_ (.A(_0593_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__clkbuf_8 _1453_ (.A(_0601_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1454_ (.A0(net416),
    .A1(_0592_),
    .S(_0000_),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _1455_ (.A(_0602_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _1456_ (.A(_0590_),
    .Y(_0284_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(net264),
    .A1(net191),
    .S(_0591_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(net415),
    .A1(_0603_),
    .S(_0000_),
    .X(_0604_));
 sky130_fd_sc_hd__clkbuf_1 _1459_ (.A(_0604_),
    .X(_0415_));
 sky130_fd_sc_hd__inv_2 _1460_ (.A(_0590_),
    .Y(_0282_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(net262),
    .A1(net189),
    .S(_0591_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(net413),
    .A1(_0605_),
    .S(_0000_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_1 _1463_ (.A(_0606_),
    .X(_0414_));
 sky130_fd_sc_hd__inv_2 _1464_ (.A(_0590_),
    .Y(_0280_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(net261),
    .A1(net188),
    .S(_0591_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _1466_ (.A0(net412),
    .A1(_0607_),
    .S(_0000_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _1467_ (.A(_0608_),
    .X(_0413_));
 sky130_fd_sc_hd__inv_2 _1468_ (.A(_0590_),
    .Y(_0278_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(net260),
    .A1(net187),
    .S(_0591_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _1470_ (.A0(net411),
    .A1(_0609_),
    .S(_0000_),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_1 _1471_ (.A(_0610_),
    .X(_0412_));
 sky130_fd_sc_hd__inv_2 _1472_ (.A(_0590_),
    .Y(_0276_));
 sky130_fd_sc_hd__mux2_1 _1473_ (.A0(net259),
    .A1(net186),
    .S(_0591_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(net410),
    .A1(_0611_),
    .S(_0000_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_1 _1475_ (.A(_0612_),
    .X(_0411_));
 sky130_fd_sc_hd__inv_2 _1476_ (.A(_0590_),
    .Y(_0274_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(net258),
    .A1(net185),
    .S(_0591_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(net409),
    .A1(_0613_),
    .S(_0000_),
    .X(_0614_));
 sky130_fd_sc_hd__clkbuf_1 _1479_ (.A(_0614_),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _1480_ (.A(_0590_),
    .Y(_0272_));
 sky130_fd_sc_hd__mux2_1 _1481_ (.A0(net257),
    .A1(net184),
    .S(_0591_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(net408),
    .A1(_0615_),
    .S(_0000_),
    .X(_0616_));
 sky130_fd_sc_hd__clkbuf_1 _1483_ (.A(_0616_),
    .X(_0409_));
 sky130_fd_sc_hd__inv_2 _1484_ (.A(_0590_),
    .Y(_0270_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(net256),
    .A1(net183),
    .S(_0591_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(net407),
    .A1(_0617_),
    .S(_0000_),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_1 _1487_ (.A(_0618_),
    .X(_0408_));
 sky130_fd_sc_hd__inv_2 _1488_ (.A(_0590_),
    .Y(_0268_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(net255),
    .A1(net182),
    .S(_0591_),
    .X(_0619_));
 sky130_fd_sc_hd__buf_4 _1490_ (.A(_0601_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _1491_ (.A0(net406),
    .A1(_0619_),
    .S(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_0621_),
    .X(_0407_));
 sky130_fd_sc_hd__buf_6 _1493_ (.A(_0589_),
    .X(_0622_));
 sky130_fd_sc_hd__inv_2 _1494_ (.A(_0622_),
    .Y(_0266_));
 sky130_fd_sc_hd__buf_4 _1495_ (.A(net205),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(net254),
    .A1(net181),
    .S(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(net405),
    .A1(_0624_),
    .S(_0620_),
    .X(_0625_));
 sky130_fd_sc_hd__clkbuf_1 _1498_ (.A(_0625_),
    .X(_0406_));
 sky130_fd_sc_hd__inv_2 _1499_ (.A(_0622_),
    .Y(_0264_));
 sky130_fd_sc_hd__mux2_1 _1500_ (.A0(net253),
    .A1(net180),
    .S(_0623_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _1501_ (.A0(net404),
    .A1(_0626_),
    .S(_0620_),
    .X(_0627_));
 sky130_fd_sc_hd__clkbuf_1 _1502_ (.A(_0627_),
    .X(_0405_));
 sky130_fd_sc_hd__inv_2 _1503_ (.A(_0622_),
    .Y(_0262_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(net251),
    .A1(net178),
    .S(_0623_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(net402),
    .A1(_0628_),
    .S(_0620_),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_1 _1506_ (.A(_0629_),
    .X(_0404_));
 sky130_fd_sc_hd__inv_2 _1507_ (.A(_0622_),
    .Y(_0260_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(net250),
    .A1(net177),
    .S(_0623_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _1509_ (.A0(net401),
    .A1(_0630_),
    .S(_0620_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _1510_ (.A(_0631_),
    .X(_0403_));
 sky130_fd_sc_hd__inv_2 _1511_ (.A(_0622_),
    .Y(_0258_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(net249),
    .A1(net176),
    .S(_0623_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(net400),
    .A1(_0632_),
    .S(_0620_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1514_ (.A(_0633_),
    .X(_0402_));
 sky130_fd_sc_hd__inv_2 _1515_ (.A(_0622_),
    .Y(_0256_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(net248),
    .A1(net175),
    .S(_0623_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(net399),
    .A1(_0634_),
    .S(_0620_),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _1518_ (.A(_0635_),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _1519_ (.A(_0622_),
    .Y(_0254_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(net247),
    .A1(net174),
    .S(_0623_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _1521_ (.A0(net398),
    .A1(_0636_),
    .S(_0620_),
    .X(_0637_));
 sky130_fd_sc_hd__clkbuf_1 _1522_ (.A(_0637_),
    .X(_0400_));
 sky130_fd_sc_hd__inv_2 _1523_ (.A(_0622_),
    .Y(_0252_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(net246),
    .A1(net173),
    .S(_0623_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(net397),
    .A1(_0638_),
    .S(_0620_),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_0639_),
    .X(_0399_));
 sky130_fd_sc_hd__inv_2 _1527_ (.A(_0622_),
    .Y(_0250_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(net245),
    .A1(net172),
    .S(_0623_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(net396),
    .A1(_0640_),
    .S(_0620_),
    .X(_0641_));
 sky130_fd_sc_hd__clkbuf_1 _1530_ (.A(_0641_),
    .X(_0398_));
 sky130_fd_sc_hd__inv_2 _1531_ (.A(_0622_),
    .Y(_0248_));
 sky130_fd_sc_hd__mux2_1 _1532_ (.A0(net244),
    .A1(net171),
    .S(_0623_),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_8 _1533_ (.A(_0601_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(net395),
    .A1(_0642_),
    .S(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__clkbuf_1 _1535_ (.A(_0644_),
    .X(_0397_));
 sky130_fd_sc_hd__buf_6 _1536_ (.A(_0589_),
    .X(_0645_));
 sky130_fd_sc_hd__inv_2 _1537_ (.A(_0645_),
    .Y(_0246_));
 sky130_fd_sc_hd__buf_4 _1538_ (.A(net205),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _1539_ (.A0(net243),
    .A1(net170),
    .S(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(net394),
    .A1(_0647_),
    .S(_0643_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_1 _1541_ (.A(_0648_),
    .X(_0396_));
 sky130_fd_sc_hd__inv_2 _1542_ (.A(_0645_),
    .Y(_0244_));
 sky130_fd_sc_hd__mux2_1 _1543_ (.A0(net242),
    .A1(net169),
    .S(_0646_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(net393),
    .A1(_0649_),
    .S(_0643_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_1 _1545_ (.A(_0650_),
    .X(_0395_));
 sky130_fd_sc_hd__inv_2 _1546_ (.A(_0645_),
    .Y(_0242_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(net272),
    .A1(net210),
    .S(_0646_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(net423),
    .A1(_0651_),
    .S(_0643_),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_1 _1549_ (.A(_0652_),
    .X(_0394_));
 sky130_fd_sc_hd__inv_2 _1550_ (.A(_0645_),
    .Y(_0240_));
 sky130_fd_sc_hd__mux2_1 _1551_ (.A0(net271),
    .A1(net209),
    .S(_0646_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(net422),
    .A1(_0653_),
    .S(_0643_),
    .X(_0654_));
 sky130_fd_sc_hd__clkbuf_1 _1553_ (.A(_0654_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _1554_ (.A(_0645_),
    .Y(_0238_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(net270),
    .A1(net208),
    .S(_0646_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(net421),
    .A1(_0655_),
    .S(_0643_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _1557_ (.A(_0656_),
    .X(_0392_));
 sky130_fd_sc_hd__inv_2 _1558_ (.A(_0645_),
    .Y(_0236_));
 sky130_fd_sc_hd__mux2_1 _1559_ (.A0(net269),
    .A1(net207),
    .S(_0646_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(net420),
    .A1(_0657_),
    .S(_0643_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _1561_ (.A(_0658_),
    .X(_0391_));
 sky130_fd_sc_hd__inv_2 _1562_ (.A(_0645_),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(net268),
    .A1(net204),
    .S(_0646_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net419),
    .A1(_0659_),
    .S(_0643_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _1565_ (.A(_0660_),
    .X(_0390_));
 sky130_fd_sc_hd__inv_2 _1566_ (.A(_0645_),
    .Y(_0232_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(net267),
    .A1(net203),
    .S(_0646_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(net418),
    .A1(_0661_),
    .S(_0643_),
    .X(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _1569_ (.A(_0662_),
    .X(_0389_));
 sky130_fd_sc_hd__inv_2 _1570_ (.A(_0645_),
    .Y(_0230_));
 sky130_fd_sc_hd__mux2_1 _1571_ (.A0(net266),
    .A1(net201),
    .S(_0646_),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(net417),
    .A1(_0663_),
    .S(_0643_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_1 _1573_ (.A(_0664_),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _1574_ (.A(_0645_),
    .Y(_0228_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(net263),
    .A1(net190),
    .S(_0646_),
    .X(_0665_));
 sky130_fd_sc_hd__buf_4 _1576_ (.A(_0601_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(net414),
    .A1(_0665_),
    .S(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_1 _1578_ (.A(_0667_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_6 _1579_ (.A(_0589_),
    .X(_0668_));
 sky130_fd_sc_hd__inv_2 _1580_ (.A(_0668_),
    .Y(_0226_));
 sky130_fd_sc_hd__buf_4 _1581_ (.A(net205),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(net252),
    .A1(net179),
    .S(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(net403),
    .A1(_0670_),
    .S(_0666_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _1584_ (.A(_0671_),
    .X(_0386_));
 sky130_fd_sc_hd__inv_2 _1585_ (.A(_0668_),
    .Y(_0224_));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(net241),
    .A1(net168),
    .S(_0669_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(net392),
    .A1(_0672_),
    .S(_0666_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _1588_ (.A(_0673_),
    .X(_0385_));
 sky130_fd_sc_hd__inv_2 _1589_ (.A(_0668_),
    .Y(_0222_));
 sky130_fd_sc_hd__mux2_1 _1590_ (.A0(net213),
    .A1(net202),
    .S(_0669_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _1591_ (.A0(net390),
    .A1(_0674_),
    .S(_0666_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _1592_ (.A(_0675_),
    .X(_0384_));
 sky130_fd_sc_hd__inv_2 _1593_ (.A(_0668_),
    .Y(_0220_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(net239),
    .A1(net200),
    .S(_0669_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(net389),
    .A1(_0676_),
    .S(_0666_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _1596_ (.A(_0677_),
    .X(_0383_));
 sky130_fd_sc_hd__inv_2 _1597_ (.A(_0668_),
    .Y(_0218_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(net238),
    .A1(net199),
    .S(_0669_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(net388),
    .A1(_0678_),
    .S(_0666_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_1 _1600_ (.A(_0679_),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _1601_ (.A(_0668_),
    .Y(_0216_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(net237),
    .A1(net198),
    .S(_0669_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(net387),
    .A1(_0680_),
    .S(_0666_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_1 _1604_ (.A(_0681_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _1605_ (.A(_0668_),
    .Y(_0214_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(net236),
    .A1(net197),
    .S(_0669_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(net386),
    .A1(_0682_),
    .S(_0666_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _1608_ (.A(_0683_),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _1609_ (.A(_0668_),
    .Y(_0212_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(net235),
    .A1(net196),
    .S(_0669_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _1611_ (.A0(net385),
    .A1(_0684_),
    .S(_0666_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _1612_ (.A(_0685_),
    .X(_0379_));
 sky130_fd_sc_hd__inv_2 _1613_ (.A(_0668_),
    .Y(_0210_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(net234),
    .A1(net195),
    .S(_0669_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(net384),
    .A1(_0686_),
    .S(_0666_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _1616_ (.A(_0687_),
    .X(_0378_));
 sky130_fd_sc_hd__inv_2 _1617_ (.A(_0668_),
    .Y(_0208_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(net233),
    .A1(net194),
    .S(_0669_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(net383),
    .A1(_0688_),
    .S(_0601_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _1620_ (.A(_0689_),
    .X(_0377_));
 sky130_fd_sc_hd__buf_12 _1621_ (.A(_0589_),
    .X(_0690_));
 sky130_fd_sc_hd__inv_2 _1622_ (.A(_0690_),
    .Y(_0206_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(net230),
    .A1(net193),
    .S(net205),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(prog_h_addr0),
    .A1(_0691_),
    .S(_0601_),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _1625_ (.A(_0692_),
    .X(_0376_));
 sky130_fd_sc_hd__inv_2 _1626_ (.A(_0690_),
    .Y(_0204_));
 sky130_fd_sc_hd__or4bb_1 _1627_ (.A(net219),
    .B(net212),
    .C_N(net230),
    .D_N(net233),
    .X(_0693_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0594_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__and4b_1 _1629_ (.A_N(net214),
    .B(net213),
    .C(net238),
    .D(net239),
    .X(_0695_));
 sky130_fd_sc_hd__and3_1 _1630_ (.A(net234),
    .B(net237),
    .C(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _1631_ (.A(net235),
    .B(net236),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_1 _1632_ (.A(_0599_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a31o_1 _1633_ (.A1(_0694_),
    .A2(_0696_),
    .A3(_0698_),
    .B1(net206),
    .X(_0699_));
 sky130_fd_sc_hd__a21o_1 _1634_ (.A1(_0593_),
    .A2(_0699_),
    .B1(net602),
    .X(_0375_));
 sky130_fd_sc_hd__inv_2 _1635_ (.A(_0690_),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _1636_ (.A(_0690_),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1637_ (.A(_0690_),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1638_ (.A(_0690_),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1639_ (.A(_0690_),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1640_ (.A(_0690_),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1641_ (.A(_0690_),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1642_ (.A(_0690_),
    .Y(_0156_));
 sky130_fd_sc_hd__buf_6 _1643_ (.A(_0589_),
    .X(_0700_));
 sky130_fd_sc_hd__inv_2 _1644_ (.A(_0700_),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1645_ (.A(_0700_),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(_0700_),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(_0700_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1648_ (.A(_0700_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1649_ (.A(_0700_),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1650_ (.A(_0700_),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1651_ (.A(_0700_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1652_ (.A(_0700_),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1653_ (.A(_0700_),
    .Y(_0136_));
 sky130_fd_sc_hd__buf_6 _1654_ (.A(_0589_),
    .X(_0701_));
 sky130_fd_sc_hd__inv_2 _1655_ (.A(_0701_),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1656_ (.A(_0701_),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1657_ (.A(_0701_),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1658_ (.A(_0701_),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1659_ (.A(_0701_),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1660_ (.A(_0701_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1661_ (.A(_0701_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1662_ (.A(_0701_),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1663_ (.A(_0701_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1664_ (.A(_0701_),
    .Y(_0116_));
 sky130_fd_sc_hd__buf_6 _1665_ (.A(_0589_),
    .X(_0702_));
 sky130_fd_sc_hd__inv_2 _1666_ (.A(_0702_),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1667_ (.A(_0702_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1668_ (.A(_0702_),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1669_ (.A(_0702_),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1670_ (.A(_0702_),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1671_ (.A(_0702_),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1672_ (.A(_0702_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1673_ (.A(_0702_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1674_ (.A(_0702_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1675_ (.A(_0702_),
    .Y(_0096_));
 sky130_fd_sc_hd__buf_6 _1676_ (.A(net211),
    .X(_0703_));
 sky130_fd_sc_hd__inv_2 _1677_ (.A(_0703_),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1678_ (.A(_0703_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1679_ (.A(_0703_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1680_ (.A(_0703_),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1681_ (.A(_0703_),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1682_ (.A(_0703_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1683_ (.A(_0703_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1684_ (.A(_0703_),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1685_ (.A(_0703_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1686_ (.A(_0703_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1687_ (.A(_0589_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1688_ (.A(_0589_),
    .Y(_0072_));
 sky130_fd_sc_hd__and2_1 _1689_ (.A(\i_ca.ca_wr_et_const ),
    .B(\i_ca.ca_ready ),
    .X(_0704_));
 sky130_fd_sc_hd__or2b_4 _1690_ (.A(\i_ca.ca_wr_com_const ),
    .B_N(\i_ca.ca_wr_fsm_state[9] ),
    .X(_0705_));
 sky130_fd_sc_hd__or2_1 _1691_ (.A(_0704_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__inv_2 _1692_ (.A(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21a_1 _1693_ (.A1(\i_ca.ca_wr_fsm_state[14] ),
    .A2(_0707_),
    .B1(\i_ca.ca_wr_sync_update ),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_8 _1694_ (.A(\i_ca.ca_wr_add_start_marker ),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_2 _1695_ (.A0(\i_ca.ca_insert_lesser_high ),
    .A1(\i_ca.ca_insert_lesser_low ),
    .S(\i_ca.ca_insert_equal_high ),
    .X(_0709_));
 sky130_fd_sc_hd__and4_1 _1696_ (.A(_0708_),
    .B(\i_ca.ca_compare_check ),
    .C(\i_ca.ca_wr_fsm_state[16] ),
    .D(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__and2b_2 _1697_ (.A_N(\i_ca.ca_wr_douta[32] ),
    .B(\i_ca.ca_wr_fsm_state[7] ),
    .X(_0711_));
 sky130_fd_sc_hd__a2111o_1 _1698_ (.A1(\i_ca.ca_wr_fsm_state[1] ),
    .A2(\i_ca.ca_wr_douta[32] ),
    .B1(\i_ca.ca_wr_fsm_state[4] ),
    .C1(_0710_),
    .D1(_0711_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_2 _1699_ (.A(\i_ca.ca_wr_add[0] ),
    .B(\i_ca.ca_wr_add[1] ),
    .C(\i_ca.ca_wr_add[2] ),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _1700_ (.A(\i_ca.ca_wr_add[3] ),
    .B(\i_ca.ca_wr_add[4] ),
    .C(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__and2_1 _1701_ (.A(\i_ca.ca_wr_add[5] ),
    .B(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__or4b_2 _1702_ (.A(\i_ca.ca_wr_add[7] ),
    .B(\i_ca.ca_wr_add[6] ),
    .C(\i_ca.ca_wr_add[8] ),
    .D_N(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__inv_2 _1703_ (.A(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nor2_1 _1704_ (.A(\i_ca.ca_wr_sync_update ),
    .B(_0706_),
    .Y(_0717_));
 sky130_fd_sc_hd__inv_2 _1705_ (.A(\i_ca.ca_wr_sync_update ),
    .Y(_0718_));
 sky130_fd_sc_hd__buf_4 _1706_ (.A(\i_ca.ca_wr_fsm_state[9] ),
    .X(_0719_));
 sky130_fd_sc_hd__buf_4 _1707_ (.A(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__and2b_1 _1708_ (.A_N(\i_ca.ca_wr_douta[32] ),
    .B(\i_ca.ca_wr_fsm_state[1] ),
    .X(_0721_));
 sky130_fd_sc_hd__a221o_1 _1709_ (.A1(\i_ca.ca_wr_fsm_state[14] ),
    .A2(_0718_),
    .B1(\i_ca.ca_wr_com_const ),
    .B2(_0720_),
    .C1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__a211o_1 _1710_ (.A1(\i_ca.ca_wr_fsm_state[0] ),
    .A2(_0716_),
    .B1(_0717_),
    .C1(_0722_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _1711_ (.A(\i_ca.ca_update_rd_add ),
    .Y(_0723_));
 sky130_fd_sc_hd__inv_2 _1712_ (.A(\i_ca.ca_match_block_ack ),
    .Y(_0724_));
 sky130_fd_sc_hd__and2_1 _1713_ (.A(_0723_),
    .B(\i_ca.ca_rd_fsm_state[2] ),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_2 _1714_ (.A(_0725_),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _1715_ (.A1(\i_ca.ca_rd_fsm_state[7] ),
    .A2(_0723_),
    .B1(_0724_),
    .B2(_0034_),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _1716_ (.A(\i_ca.ca_match_ack_meta ),
    .Y(_0726_));
 sky130_fd_sc_hd__inv_2 _1717_ (.A(\i_ca.ca_match_req ),
    .Y(_0727_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(\i_ca.ca_match_hs_state[0] ),
    .B(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__a21o_1 _1719_ (.A1(\i_ca.ca_match_hs_state[1] ),
    .A2(_0726_),
    .B1(_0728_),
    .X(_0016_));
 sky130_fd_sc_hd__inv_2 _1720_ (.A(\i_ca.ca_insert_time[11] ),
    .Y(_0729_));
 sky130_fd_sc_hd__inv_2 _1721_ (.A(\i_ca.ca_insert_time[12] ),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _1722_ (.A(\i_ca.ca_insert_time[13] ),
    .Y(_0731_));
 sky130_fd_sc_hd__or2_1 _1723_ (.A(\i_ca.ca_wr_douta[13] ),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__o221a_1 _1724_ (.A1(\i_ca.ca_wr_douta[11] ),
    .A2(_0729_),
    .B1(\i_ca.ca_wr_douta[12] ),
    .B2(_0730_),
    .C1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__inv_2 _1725_ (.A(\i_ca.ca_insert_time[14] ),
    .Y(_0734_));
 sky130_fd_sc_hd__inv_2 _1726_ (.A(\i_ca.ca_insert_time[15] ),
    .Y(_0735_));
 sky130_fd_sc_hd__o22a_1 _1727_ (.A1(\i_ca.ca_wr_douta[14] ),
    .A2(_0734_),
    .B1(\i_ca.ca_wr_douta[15] ),
    .B2(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__inv_2 _1728_ (.A(\i_ca.ca_wr_douta[18] ),
    .Y(_0737_));
 sky130_fd_sc_hd__inv_2 _1729_ (.A(\i_ca.ca_insert_time[17] ),
    .Y(_0738_));
 sky130_fd_sc_hd__o2bb2a_1 _1730_ (.A1_N(_0737_),
    .A2_N(\i_ca.ca_insert_time[18] ),
    .B1(\i_ca.ca_wr_douta[17] ),
    .B2(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__inv_2 _1731_ (.A(\i_ca.ca_wr_douta[16] ),
    .Y(_0740_));
 sky130_fd_sc_hd__o2bb2a_1 _1732_ (.A1_N(_0735_),
    .A2_N(\i_ca.ca_wr_douta[15] ),
    .B1(\i_ca.ca_insert_time[16] ),
    .B2(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__and3_1 _1733_ (.A(_0736_),
    .B(_0739_),
    .C(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__inv_2 _1734_ (.A(\i_ca.ca_wr_douta[20] ),
    .Y(_0743_));
 sky130_fd_sc_hd__inv_2 _1735_ (.A(\i_ca.ca_wr_douta[21] ),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_1 _1736_ (.A(\i_ca.ca_insert_time[22] ),
    .B(\i_ca.ca_wr_douta[22] ),
    .Y(_0745_));
 sky130_fd_sc_hd__o21a_1 _1737_ (.A1(\i_ca.ca_insert_time[21] ),
    .A2(_0744_),
    .B1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a21bo_1 _1738_ (.A1(\i_ca.ca_insert_time[21] ),
    .A2(_0744_),
    .B1_N(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__a21o_1 _1739_ (.A1(_0743_),
    .A2(\i_ca.ca_insert_time[20] ),
    .B1(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__inv_2 _1740_ (.A(\i_ca.ca_wr_douta[19] ),
    .Y(_0749_));
 sky130_fd_sc_hd__and2_1 _1741_ (.A(_0749_),
    .B(\i_ca.ca_insert_time[19] ),
    .X(_0750_));
 sky130_fd_sc_hd__a22o_1 _1742_ (.A1(\i_ca.ca_wr_douta[12] ),
    .A2(_0730_),
    .B1(\i_ca.ca_wr_douta[13] ),
    .B2(_0731_),
    .X(_0751_));
 sky130_fd_sc_hd__nand2_1 _1743_ (.A(\i_ca.ca_wr_douta[11] ),
    .B(_0729_),
    .Y(_0752_));
 sky130_fd_sc_hd__inv_2 _1744_ (.A(\i_ca.ca_wr_douta[14] ),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(_0740_),
    .B(\i_ca.ca_insert_time[16] ),
    .Y(_0754_));
 sky130_fd_sc_hd__o221a_1 _1746_ (.A1(_0753_),
    .A2(\i_ca.ca_insert_time[14] ),
    .B1(_0737_),
    .B2(\i_ca.ca_insert_time[18] ),
    .C1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__nand2_1 _1747_ (.A(\i_ca.ca_wr_douta[17] ),
    .B(_0738_),
    .Y(_0756_));
 sky130_fd_sc_hd__and4b_1 _1748_ (.A_N(_0751_),
    .B(_0752_),
    .C(_0755_),
    .D(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__o22a_1 _1749_ (.A1(_0743_),
    .A2(\i_ca.ca_insert_time[20] ),
    .B1(_0749_),
    .B2(\i_ca.ca_insert_time[19] ),
    .X(_0758_));
 sky130_fd_sc_hd__and4bb_1 _1750_ (.A_N(_0748_),
    .B_N(_0750_),
    .C(_0757_),
    .D(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__and3_1 _1751_ (.A(_0733_),
    .B(_0742_),
    .C(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__clkbuf_1 _1752_ (.A(_0760_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _1753_ (.A(\i_ca.ca_wr_fsm_state[7] ),
    .B(\i_ca.ca_wr_douta[32] ),
    .X(_0761_));
 sky130_fd_sc_hd__buf_4 _1754_ (.A(_0761_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1755_ (.A(\i_ca.ca_match_hs_state[0] ),
    .B(\i_ca.ca_match_req ),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_1 _1756_ (.A(_0762_),
    .X(_0005_));
 sky130_fd_sc_hd__a21o_1 _1757_ (.A1(\i_ca.ca_match_hs_state[2] ),
    .A2(_0726_),
    .B1(_0005_),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_1 _1758_ (.A1(\i_ca.ca_wr_sync_update_done ),
    .A2(\i_ca.ca_rd_fsm_state[1] ),
    .B1(\i_ca.ca_rd_fsm_state[8] ),
    .Y(_0763_));
 sky130_fd_sc_hd__nor2_1 _1759_ (.A(\i_ca.ca_update_rd_add ),
    .B(_0763_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1760_ (.A(\i_ca.ca_wr_fsm_state[0] ),
    .Y(_0764_));
 sky130_fd_sc_hd__nor2_1 _1761_ (.A(_0764_),
    .B(_0716_),
    .Y(_0010_));
 sky130_fd_sc_hd__or2_1 _1762_ (.A(\i_ca.ca_wr_fsm_state[11] ),
    .B(\i_ca.ca_wr_fsm_state[2] ),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_1 _1763_ (.A(_0765_),
    .X(_0026_));
 sky130_fd_sc_hd__and2b_1 _1764_ (.A_N(\i_ca.ca_ready ),
    .B(\i_ca.hs_state_write_const[1] ),
    .X(_0766_));
 sky130_fd_sc_hd__or2_1 _1765_ (.A(\i_ca.hs_state_write_const[2] ),
    .B(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__clkbuf_1 _1766_ (.A(_0767_),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_4 _1767_ (.A(\i_ca.ca_compare_check ),
    .B(_0709_),
    .Y(_0768_));
 sky130_fd_sc_hd__and3_1 _1768_ (.A(\i_ca.ca_end_of_wr_list ),
    .B(\i_ca.ca_wr_fsm_state[16] ),
    .C(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__or2_1 _1769_ (.A(\i_ca.ca_wr_fsm_state[15] ),
    .B(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__buf_4 _1770_ (.A(_0770_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _1771_ (.A1(\i_ca.ca_ready ),
    .A2(\i_ca.hs_state_write_const[1] ),
    .B1(\i_ca.ca_dbus_valid_meta ),
    .B2(\i_ca.hs_state_write_const[3] ),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_1 _1772_ (.A(\i_ca.ca_wr_sync_update_done ),
    .B(\i_ca.ca_update_rd_add ),
    .Y(_0771_));
 sky130_fd_sc_hd__a22o_1 _1773_ (.A1(\i_ca.ca_match_block_ack ),
    .A2(_0034_),
    .B1(_0771_),
    .B2(\i_ca.ca_rd_fsm_state[6] ),
    .X(_0022_));
 sky130_fd_sc_hd__inv_2 _1774_ (.A(\i_ca.ca_rd_fsm_state[5] ),
    .Y(_0772_));
 sky130_fd_sc_hd__nor2_4 _1775_ (.A(\i_ca.ca_update_rd_add ),
    .B(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _1776_ (.A(\i_ca.ca_wr_add_start_marker ),
    .Y(_0774_));
 sky130_fd_sc_hd__and3_1 _1777_ (.A(\i_ca.ca_time_diff[21] ),
    .B(\i_ca.ca_time_diff[20] ),
    .C(\i_ca.ca_time_diff[22] ),
    .X(_0775_));
 sky130_fd_sc_hd__and4_1 _1778_ (.A(\i_ca.ca_time_diff[17] ),
    .B(\i_ca.ca_time_diff[16] ),
    .C(\i_ca.ca_time_diff[19] ),
    .D(\i_ca.ca_time_diff[18] ),
    .X(_0776_));
 sky130_fd_sc_hd__and4_1 _1779_ (.A(\i_ca.ca_time_diff[13] ),
    .B(\i_ca.ca_time_diff[12] ),
    .C(\i_ca.ca_time_diff[15] ),
    .D(\i_ca.ca_time_diff[14] ),
    .X(_0777_));
 sky130_fd_sc_hd__inv_2 _1780_ (.A(\i_ca.ca_match_check ),
    .Y(_0778_));
 sky130_fd_sc_hd__a31o_1 _1781_ (.A1(_0775_),
    .A2(_0776_),
    .A3(_0777_),
    .B1(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__nand3_2 _1782_ (.A(_0774_),
    .B(\i_ca.ca_rd_doutb_32 ),
    .C(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__and3_1 _1783_ (.A(\i_ca.ca_ready ),
    .B(_0723_),
    .C(\i_ca.ca_rd_fsm_state[0] ),
    .X(_0781_));
 sky130_fd_sc_hd__a221o_1 _1784_ (.A1(net874),
    .A2(_0771_),
    .B1(_0773_),
    .B2(_0780_),
    .C1(_0781_),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _1785_ (.A1(\i_ca.ca_wr_sync_update_done ),
    .A2(\i_ca.ca_rd_fsm_state[6] ),
    .B1(\i_ca.ca_update_rd_add ),
    .X(_0020_));
 sky130_fd_sc_hd__or4_1 _1786_ (.A(\i_ca.ca_rd_doutb[28] ),
    .B(\i_ca.ca_rd_doutb[27] ),
    .C(\i_ca.ca_rd_doutb[30] ),
    .D(\i_ca.ca_rd_doutb[29] ),
    .X(_0782_));
 sky130_fd_sc_hd__or4_1 _1787_ (.A(\i_ca.ca_rd_doutb[24] ),
    .B(\i_ca.ca_rd_doutb[23] ),
    .C(\i_ca.ca_rd_doutb[26] ),
    .D(\i_ca.ca_rd_doutb[25] ),
    .X(_0783_));
 sky130_fd_sc_hd__or2_1 _1788_ (.A(_0782_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(_0784_),
    .X(_0035_));
 sky130_fd_sc_hd__or4_1 _1790_ (.A(\i_ca.ca_wr_douta[28] ),
    .B(\i_ca.ca_wr_douta[27] ),
    .C(\i_ca.ca_wr_douta[30] ),
    .D(\i_ca.ca_wr_douta[29] ),
    .X(_0785_));
 sky130_fd_sc_hd__or4_1 _1791_ (.A(\i_ca.ca_wr_douta[24] ),
    .B(\i_ca.ca_wr_douta[23] ),
    .C(\i_ca.ca_wr_douta[26] ),
    .D(\i_ca.ca_wr_douta[25] ),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_1 _1792_ (.A(_0785_),
    .B(_0786_),
    .Y(_0031_));
 sky130_fd_sc_hd__buf_4 _1793_ (.A(_0769_),
    .X(_0787_));
 sky130_fd_sc_hd__nand2_4 _1794_ (.A(\i_ca.ca_wr_et_const ),
    .B(\i_ca.ca_ready ),
    .Y(_0788_));
 sky130_fd_sc_hd__a21o_1 _1795_ (.A1(\i_ca.ca_wr_sync_update ),
    .A2(_0788_),
    .B1(\i_ca.ca_wr_com_const ),
    .X(_0789_));
 sky130_fd_sc_hd__buf_4 _1796_ (.A(\i_ca.ca_wr_fsm_state[3] ),
    .X(_0790_));
 sky130_fd_sc_hd__or4_1 _1797_ (.A(\i_ca.ca_wr_fsm_state[0] ),
    .B(_0790_),
    .C(\i_ca.ca_wr_fsm_state[15] ),
    .D(_0711_),
    .X(_0791_));
 sky130_fd_sc_hd__a211o_1 _1798_ (.A1(_0719_),
    .A2(_0789_),
    .B1(_0791_),
    .C1(\i_ca.ca_wr_fsm_state[4] ),
    .X(_0792_));
 sky130_fd_sc_hd__or3_2 _1799_ (.A(_0710_),
    .B(_0787_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__clkbuf_1 _1800_ (.A(_0793_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_4 _1801_ (.A(prog_h_addr0),
    .B(prog_wea),
    .Y(net424));
 sky130_fd_sc_hd__or2b_1 _1802_ (.A(prog_h_addr0),
    .B_N(prog_wea),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_1 _1803_ (.A(_0794_),
    .X(net466));
 sky130_fd_sc_hd__inv_2 _1804_ (.A(\i_ca.ca_insert_time[10] ),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_2 _1805_ (.A(\i_ca.ca_insert_time[8] ),
    .Y(_0796_));
 sky130_fd_sc_hd__nor2_1 _1806_ (.A(_0796_),
    .B(\i_ca.ca_wr_douta[8] ),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _1807_ (.A(\i_ca.ca_insert_time[9] ),
    .Y(_0798_));
 sky130_fd_sc_hd__a22o_1 _1808_ (.A1(_0796_),
    .A2(\i_ca.ca_wr_douta[8] ),
    .B1(_0798_),
    .B2(\i_ca.ca_wr_douta[9] ),
    .X(_0799_));
 sky130_fd_sc_hd__or2_1 _1809_ (.A(_0798_),
    .B(\i_ca.ca_wr_douta[9] ),
    .X(_0800_));
 sky130_fd_sc_hd__or3b_1 _1810_ (.A(_0797_),
    .B(_0799_),
    .C_N(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__inv_2 _1811_ (.A(\i_ca.ca_insert_time[6] ),
    .Y(_0802_));
 sky130_fd_sc_hd__inv_2 _1812_ (.A(\i_ca.ca_insert_time[7] ),
    .Y(_0803_));
 sky130_fd_sc_hd__a22o_1 _1813_ (.A1(_0802_),
    .A2(\i_ca.ca_wr_douta[6] ),
    .B1(_0803_),
    .B2(\i_ca.ca_wr_douta[7] ),
    .X(_0804_));
 sky130_fd_sc_hd__or2_1 _1814_ (.A(_0803_),
    .B(\i_ca.ca_wr_douta[7] ),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _1815_ (.A(_0802_),
    .B(\i_ca.ca_wr_douta[6] ),
    .Y(_0806_));
 sky130_fd_sc_hd__or3b_1 _1816_ (.A(_0806_),
    .B(_0804_),
    .C_N(_0805_),
    .X(_0807_));
 sky130_fd_sc_hd__inv_2 _1817_ (.A(\i_ca.ca_wr_douta[2] ),
    .Y(_0808_));
 sky130_fd_sc_hd__inv_2 _1818_ (.A(\i_ca.ca_wr_douta[3] ),
    .Y(_0809_));
 sky130_fd_sc_hd__inv_2 _1819_ (.A(\i_ca.ca_insert_time[1] ),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _1820_ (.A(_0810_),
    .B(\i_ca.ca_wr_douta[1] ),
    .Y(_0811_));
 sky130_fd_sc_hd__inv_2 _1821_ (.A(\i_ca.ca_insert_time[0] ),
    .Y(_0812_));
 sky130_fd_sc_hd__o22a_1 _1822_ (.A1(_0812_),
    .A2(\i_ca.ca_wr_douta[0] ),
    .B1(_0810_),
    .B2(\i_ca.ca_wr_douta[1] ),
    .X(_0813_));
 sky130_fd_sc_hd__nand2_1 _1823_ (.A(_0811_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a22o_1 _1824_ (.A1(\i_ca.ca_insert_time[2] ),
    .A2(_0808_),
    .B1(_0811_),
    .B2(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__o221a_1 _1825_ (.A1(\i_ca.ca_insert_time[2] ),
    .A2(_0808_),
    .B1(\i_ca.ca_insert_time[3] ),
    .B2(_0809_),
    .C1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(\i_ca.ca_wr_douta[4] ),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(\i_ca.ca_wr_douta[5] ),
    .Y(_0818_));
 sky130_fd_sc_hd__o22a_1 _1828_ (.A1(\i_ca.ca_insert_time[4] ),
    .A2(_0817_),
    .B1(\i_ca.ca_insert_time[5] ),
    .B2(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__and2_1 _1829_ (.A(\i_ca.ca_insert_time[5] ),
    .B(_0818_),
    .X(_0820_));
 sky130_fd_sc_hd__a21oi_1 _1830_ (.A1(\i_ca.ca_insert_time[4] ),
    .A2(_0817_),
    .B1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand2_1 _1831_ (.A(_0819_),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _1832_ (.A(\i_ca.ca_insert_time[3] ),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_1 _1833_ (.A(_0823_),
    .B(\i_ca.ca_wr_douta[3] ),
    .Y(_0824_));
 sky130_fd_sc_hd__o32a_1 _1834_ (.A1(_0816_),
    .A2(_0822_),
    .A3(_0824_),
    .B1(_0820_),
    .B2(_0819_),
    .X(_0825_));
 sky130_fd_sc_hd__o2bb2a_1 _1835_ (.A1_N(_0804_),
    .A2_N(_0805_),
    .B1(_0807_),
    .B2(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__a2bb2o_1 _1836_ (.A1_N(_0801_),
    .A2_N(_0826_),
    .B1(_0799_),
    .B2(_0800_),
    .X(_0827_));
 sky130_fd_sc_hd__or4_1 _1837_ (.A(_0801_),
    .B(_0807_),
    .C(_0814_),
    .D(_0822_),
    .X(_0828_));
 sky130_fd_sc_hd__inv_2 _1838_ (.A(\i_ca.ca_insert_time[2] ),
    .Y(_0829_));
 sky130_fd_sc_hd__a221o_1 _1839_ (.A1(_0812_),
    .A2(\i_ca.ca_wr_douta[0] ),
    .B1(\i_ca.ca_insert_time[2] ),
    .B2(_0808_),
    .C1(_0824_),
    .X(_0830_));
 sky130_fd_sc_hd__a221o_1 _1840_ (.A1(_0829_),
    .A2(\i_ca.ca_wr_douta[2] ),
    .B1(_0823_),
    .B2(\i_ca.ca_wr_douta[3] ),
    .C1(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__o22a_1 _1841_ (.A1(_0795_),
    .A2(\i_ca.ca_wr_douta[10] ),
    .B1(_0828_),
    .B2(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__a22o_1 _1842_ (.A1(_0795_),
    .A2(\i_ca.ca_wr_douta[10] ),
    .B1(_0827_),
    .B2(_0832_),
    .X(_0028_));
 sky130_fd_sc_hd__or4_1 _1843_ (.A(\i_ca.ca_time_const[15] ),
    .B(\i_ca.ca_time_const[14] ),
    .C(\i_ca.ca_time_const[17] ),
    .D(\i_ca.ca_time_const[16] ),
    .X(_0833_));
 sky130_fd_sc_hd__and4b_1 _1844_ (.A_N(\i_ca.ca_time_const[22] ),
    .B(\i_ca.ca_rd_doutb[13] ),
    .C(\i_ca.ca_rd_doutb[12] ),
    .D(\i_ca.ca_rd_doutb[15] ),
    .X(_0834_));
 sky130_fd_sc_hd__or4b_1 _1845_ (.A(\i_ca.ca_time_const[19] ),
    .B(\i_ca.ca_time_const[18] ),
    .C(\i_ca.ca_time_const[21] ),
    .D_N(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__nand4_1 _1846_ (.A(\i_ca.ca_rd_doutb[18] ),
    .B(\i_ca.ca_rd_doutb[21] ),
    .C(\i_ca.ca_rd_doutb[20] ),
    .D(\i_ca.ca_rd_doutb[22] ),
    .Y(_0836_));
 sky130_fd_sc_hd__and4_1 _1847_ (.A(\i_ca.ca_rd_doutb[14] ),
    .B(\i_ca.ca_rd_doutb[17] ),
    .C(\i_ca.ca_rd_doutb[16] ),
    .D(\i_ca.ca_rd_doutb[19] ),
    .X(_0837_));
 sky130_fd_sc_hd__or4b_1 _1848_ (.A(\i_ca.ca_time_const[20] ),
    .B(_0835_),
    .C(_0836_),
    .D_N(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__or4_1 _1849_ (.A(\i_ca.ca_time_const[13] ),
    .B(\i_ca.ca_time_const[12] ),
    .C(_0833_),
    .D(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_1 _1850_ (.A(_0839_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(\i_ca.ca_wr_wea ),
    .Y(\i_ca.cubev_ca_wea ));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(\i_ca.ca_time_const[0] ),
    .Y(_0038_));
 sky130_fd_sc_hd__xor2_1 _1853_ (.A(net104),
    .B(net136),
    .X(net564));
 sky130_fd_sc_hd__xor2_1 _1854_ (.A(net115),
    .B(net147),
    .X(net575));
 sky130_fd_sc_hd__xor2_1 _1855_ (.A(net126),
    .B(net158),
    .X(net586));
 sky130_fd_sc_hd__xor2_1 _1856_ (.A(net129),
    .B(net161),
    .X(net589));
 sky130_fd_sc_hd__xor2_1 _1857_ (.A(net130),
    .B(net162),
    .X(net590));
 sky130_fd_sc_hd__xor2_1 _1858_ (.A(net131),
    .B(net163),
    .X(net591));
 sky130_fd_sc_hd__xor2_1 _1859_ (.A(net132),
    .B(net164),
    .X(net592));
 sky130_fd_sc_hd__xor2_1 _1860_ (.A(net133),
    .B(net165),
    .X(net593));
 sky130_fd_sc_hd__xor2_1 _1861_ (.A(net134),
    .B(net166),
    .X(net594));
 sky130_fd_sc_hd__xor2_1 _1862_ (.A(net135),
    .B(net167),
    .X(net595));
 sky130_fd_sc_hd__xor2_1 _1863_ (.A(net105),
    .B(net137),
    .X(net565));
 sky130_fd_sc_hd__xor2_1 _1864_ (.A(net106),
    .B(net138),
    .X(net566));
 sky130_fd_sc_hd__xor2_2 _1865_ (.A(net107),
    .B(net139),
    .X(net567));
 sky130_fd_sc_hd__xor2_1 _1866_ (.A(net108),
    .B(net140),
    .X(net568));
 sky130_fd_sc_hd__xor2_1 _1867_ (.A(net109),
    .B(net141),
    .X(net569));
 sky130_fd_sc_hd__xor2_1 _1868_ (.A(net110),
    .B(net142),
    .X(net570));
 sky130_fd_sc_hd__xor2_1 _1869_ (.A(net111),
    .B(net143),
    .X(net571));
 sky130_fd_sc_hd__xor2_1 _1870_ (.A(net112),
    .B(net144),
    .X(net572));
 sky130_fd_sc_hd__xor2_2 _1871_ (.A(net113),
    .B(net145),
    .X(net573));
 sky130_fd_sc_hd__xor2_2 _1872_ (.A(net114),
    .B(net146),
    .X(net574));
 sky130_fd_sc_hd__xor2_1 _1873_ (.A(net116),
    .B(net148),
    .X(net576));
 sky130_fd_sc_hd__xor2_1 _1874_ (.A(net117),
    .B(net149),
    .X(net577));
 sky130_fd_sc_hd__xor2_2 _1875_ (.A(net118),
    .B(net150),
    .X(net578));
 sky130_fd_sc_hd__xor2_1 _1876_ (.A(net119),
    .B(net151),
    .X(net579));
 sky130_fd_sc_hd__xor2_2 _1877_ (.A(net120),
    .B(net152),
    .X(net580));
 sky130_fd_sc_hd__xor2_2 _1878_ (.A(net121),
    .B(net153),
    .X(net581));
 sky130_fd_sc_hd__xor2_2 _1879_ (.A(net122),
    .B(net154),
    .X(net582));
 sky130_fd_sc_hd__xor2_2 _1880_ (.A(net123),
    .B(net155),
    .X(net583));
 sky130_fd_sc_hd__xor2_2 _1881_ (.A(net124),
    .B(net156),
    .X(net584));
 sky130_fd_sc_hd__xor2_2 _1882_ (.A(net125),
    .B(net157),
    .X(net585));
 sky130_fd_sc_hd__xor2_2 _1883_ (.A(net127),
    .B(net159),
    .X(net587));
 sky130_fd_sc_hd__xor2_2 _1884_ (.A(net128),
    .B(net160),
    .X(net588));
 sky130_fd_sc_hd__and3b_1 _1885_ (.A_N(\i_ca.ca_ready ),
    .B(_0723_),
    .C(\i_ca.ca_rd_fsm_state[0] ),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _1886_ (.A(_0840_),
    .X(_0006_));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(\i_ca.ca_wr_fsm_state[16] ),
    .Y(_0841_));
 sky130_fd_sc_hd__or3_4 _1888_ (.A(\i_ca.ca_wr_add_start_marker ),
    .B(_0841_),
    .C(_0768_),
    .X(_0842_));
 sky130_fd_sc_hd__inv_2 _1889_ (.A(_0842_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1890_ (.A(_0773_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(_0843_),
    .B(_0780_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21a_1 _1892_ (.A1(\i_ca.ca_match_hs_state[2] ),
    .A2(\i_ca.ca_match_hs_state[1] ),
    .B1(\i_ca.ca_match_ack_meta ),
    .X(_0004_));
 sky130_fd_sc_hd__and3_1 _1893_ (.A(\i_ca.ca_ready ),
    .B(\i_ca.hs_state_write_const[1] ),
    .C(net1),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_1 _1894_ (.A(_0844_),
    .X(_0036_));
 sky130_fd_sc_hd__nand2_8 _1895_ (.A(\i_ca.ca_ready ),
    .B(\i_ca.hs_state_write_const[1] ),
    .Y(_0845_));
 sky130_fd_sc_hd__buf_4 _1896_ (.A(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__nor2_1 _1897_ (.A(net1),
    .B(_0846_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1898_ (.A(\i_ca.ca_wr_douta[22] ),
    .Y(_0847_));
 sky130_fd_sc_hd__a221o_1 _1899_ (.A1(\i_ca.ca_wr_douta[14] ),
    .A2(_0734_),
    .B1(_0732_),
    .B2(_0751_),
    .C1(_0733_),
    .X(_0848_));
 sky130_fd_sc_hd__a21bo_1 _1900_ (.A1(_0736_),
    .A2(_0848_),
    .B1_N(_0741_),
    .X(_0849_));
 sky130_fd_sc_hd__a21bo_1 _1901_ (.A1(_0754_),
    .A2(_0849_),
    .B1_N(_0756_),
    .X(_0850_));
 sky130_fd_sc_hd__o2bb2a_1 _1902_ (.A1_N(_0850_),
    .A2_N(_0739_),
    .B1(\i_ca.ca_insert_time[18] ),
    .B2(_0737_),
    .X(_0851_));
 sky130_fd_sc_hd__o21a_1 _1903_ (.A1(_0750_),
    .A2(_0851_),
    .B1(_0758_),
    .X(_0852_));
 sky130_fd_sc_hd__o22a_1 _1904_ (.A1(\i_ca.ca_insert_time[22] ),
    .A2(_0847_),
    .B1(_0748_),
    .B2(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__a21oi_1 _1905_ (.A1(\i_ca.ca_insert_time[21] ),
    .A2(_0744_),
    .B1(_0745_),
    .Y(_0854_));
 sky130_fd_sc_hd__or2_1 _1906_ (.A(_0746_),
    .B(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__o21ai_1 _1907_ (.A1(_0029_),
    .A2(_0853_),
    .B1(_0855_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _1908_ (.A(_0747_),
    .B(_0855_),
    .Y(_0030_));
 sky130_fd_sc_hd__o21ba_1 _1909_ (.A1(\i_ca.hs_state_write_const[3] ),
    .A2(\i_ca.hs_state_write_const[0] ),
    .B1_N(\i_ca.ca_dbus_valid_meta ),
    .X(_0002_));
 sky130_fd_sc_hd__and2_1 _1910_ (.A(\i_ca.ca_dbus_valid_meta ),
    .B(\i_ca.hs_state_write_const[0] ),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_1 _1911_ (.A(_0856_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_4 _1912_ (.A(_0788_),
    .B(_0705_),
    .Y(_0857_));
 sky130_fd_sc_hd__buf_6 _1913_ (.A(_0857_),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_4 _1914_ (.A(\i_ca.ca_wr_fsm_state[16] ),
    .B(_0768_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_2 _1915_ (.A(\i_ca.ca_end_of_wr_list ),
    .B(_0858_),
    .Y(_0011_));
 sky130_fd_sc_hd__and2_1 _1916_ (.A(_0723_),
    .B(\i_ca.ca_rd_fsm_state[4] ),
    .X(_0859_));
 sky130_fd_sc_hd__clkbuf_1 _1917_ (.A(_0859_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _1918_ (.A(_0723_),
    .B(\i_ca.ca_rd_fsm_state[3] ),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_1 _1919_ (.A(_0860_),
    .X(_0008_));
 sky130_fd_sc_hd__inv_2 _1920_ (.A(\i_ca.ca_rd_doutb[7] ),
    .Y(_0861_));
 sky130_fd_sc_hd__inv_2 _1921_ (.A(\i_ca.ca_rd_doutb[6] ),
    .Y(_0862_));
 sky130_fd_sc_hd__o22a_1 _1922_ (.A1(\i_ca.ca_time_const[7] ),
    .A2(_0861_),
    .B1(\i_ca.ca_time_const[6] ),
    .B2(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__inv_2 _1923_ (.A(\i_ca.ca_rd_doutb[5] ),
    .Y(_0864_));
 sky130_fd_sc_hd__inv_2 _1924_ (.A(\i_ca.ca_rd_doutb[4] ),
    .Y(_0865_));
 sky130_fd_sc_hd__o22a_1 _1925_ (.A1(\i_ca.ca_time_const[5] ),
    .A2(_0864_),
    .B1(_0865_),
    .B2(\i_ca.ca_time_const[4] ),
    .X(_0866_));
 sky130_fd_sc_hd__inv_2 _1926_ (.A(\i_ca.ca_rd_doutb[2] ),
    .Y(_0867_));
 sky130_fd_sc_hd__or2b_1 _1927_ (.A(\i_ca.ca_time_const[1] ),
    .B_N(\i_ca.ca_rd_doutb[1] ),
    .X(_0868_));
 sky130_fd_sc_hd__and2b_1 _1928_ (.A_N(\i_ca.ca_rd_doutb[0] ),
    .B(\i_ca.ca_time_const[0] ),
    .X(_0869_));
 sky130_fd_sc_hd__and2b_1 _1929_ (.A_N(\i_ca.ca_rd_doutb[1] ),
    .B(\i_ca.ca_time_const[1] ),
    .X(_0870_));
 sky130_fd_sc_hd__a221o_1 _1930_ (.A1(\i_ca.ca_time_const[2] ),
    .A2(_0867_),
    .B1(_0868_),
    .B2(_0869_),
    .C1(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__inv_2 _1931_ (.A(\i_ca.ca_rd_doutb[3] ),
    .Y(_0872_));
 sky130_fd_sc_hd__o22a_1 _1932_ (.A1(\i_ca.ca_time_const[3] ),
    .A2(_0872_),
    .B1(\i_ca.ca_time_const[2] ),
    .B2(_0867_),
    .X(_0873_));
 sky130_fd_sc_hd__a22o_1 _1933_ (.A1(_0865_),
    .A2(\i_ca.ca_time_const[4] ),
    .B1(\i_ca.ca_time_const[3] ),
    .B2(_0872_),
    .X(_0874_));
 sky130_fd_sc_hd__a21o_1 _1934_ (.A1(_0871_),
    .A2(_0873_),
    .B1(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__a22o_1 _1935_ (.A1(\i_ca.ca_time_const[6] ),
    .A2(_0862_),
    .B1(\i_ca.ca_time_const[5] ),
    .B2(_0864_),
    .X(_0876_));
 sky130_fd_sc_hd__a21o_1 _1936_ (.A1(_0866_),
    .A2(_0875_),
    .B1(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__inv_2 _1937_ (.A(\i_ca.ca_rd_doutb[8] ),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_1 _1938_ (.A(_0878_),
    .B(\i_ca.ca_time_const[8] ),
    .Y(_0879_));
 sky130_fd_sc_hd__and2b_1 _1939_ (.A_N(\i_ca.ca_time_const[9] ),
    .B(\i_ca.ca_rd_doutb[9] ),
    .X(_0880_));
 sky130_fd_sc_hd__and2b_1 _1940_ (.A_N(\i_ca.ca_time_const[10] ),
    .B(\i_ca.ca_rd_doutb[10] ),
    .X(_0881_));
 sky130_fd_sc_hd__or3_1 _1941_ (.A(_0879_),
    .B(_0880_),
    .C(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__inv_2 _1942_ (.A(\i_ca.ca_time_const[11] ),
    .Y(_0883_));
 sky130_fd_sc_hd__and2_1 _1943_ (.A(\i_ca.ca_rd_doutb[11] ),
    .B(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__a2bb2o_1 _1944_ (.A1_N(\i_ca.ca_rd_doutb[11] ),
    .A2_N(_0883_),
    .B1(\i_ca.ca_time_const[7] ),
    .B2(_0861_),
    .X(_0885_));
 sky130_fd_sc_hd__a211o_1 _1945_ (.A1(_0878_),
    .A2(\i_ca.ca_time_const[8] ),
    .B1(_0884_),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or2b_1 _1946_ (.A(\i_ca.ca_rd_doutb[10] ),
    .B_N(\i_ca.ca_time_const[10] ),
    .X(_0887_));
 sky130_fd_sc_hd__or2b_1 _1947_ (.A(\i_ca.ca_rd_doutb[9] ),
    .B_N(\i_ca.ca_time_const[9] ),
    .X(_0888_));
 sky130_fd_sc_hd__or4bb_1 _1948_ (.A(_0882_),
    .B(_0886_),
    .C_N(_0887_),
    .D_N(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__a21o_1 _1949_ (.A1(_0863_),
    .A2(_0877_),
    .B1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__or2_1 _1950_ (.A(_0879_),
    .B(_0880_),
    .X(_0891_));
 sky130_fd_sc_hd__a311o_1 _1951_ (.A1(_0888_),
    .A2(_0887_),
    .A3(_0891_),
    .B1(_0884_),
    .C1(_0881_),
    .X(_0892_));
 sky130_fd_sc_hd__o21ai_2 _1952_ (.A1(\i_ca.ca_rd_doutb[11] ),
    .A2(_0883_),
    .B1(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__xor2_2 _1953_ (.A(\i_ca.ca_time_const[12] ),
    .B(\i_ca.ca_rd_doutb[12] ),
    .X(_0894_));
 sky130_fd_sc_hd__a21o_1 _1954_ (.A1(_0890_),
    .A2(_0893_),
    .B1(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nand3_1 _1955_ (.A(_0894_),
    .B(_0890_),
    .C(_0893_),
    .Y(_0896_));
 sky130_fd_sc_hd__and2_1 _1956_ (.A(_0895_),
    .B(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__clkbuf_1 _1957_ (.A(_0897_),
    .X(_0061_));
 sky130_fd_sc_hd__and2b_1 _1958_ (.A_N(\i_ca.ca_time_const[13] ),
    .B(\i_ca.ca_rd_doutb[13] ),
    .X(_0898_));
 sky130_fd_sc_hd__and2b_1 _1959_ (.A_N(\i_ca.ca_rd_doutb[13] ),
    .B(\i_ca.ca_time_const[13] ),
    .X(_0899_));
 sky130_fd_sc_hd__nor2_1 _1960_ (.A(_0898_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__inv_2 _1961_ (.A(\i_ca.ca_rd_doutb[12] ),
    .Y(_0901_));
 sky130_fd_sc_hd__o21a_1 _1962_ (.A1(\i_ca.ca_time_const[12] ),
    .A2(_0901_),
    .B1(_0895_),
    .X(_0902_));
 sky130_fd_sc_hd__xnor2_1 _1963_ (.A(_0900_),
    .B(_0902_),
    .Y(_0062_));
 sky130_fd_sc_hd__or2b_1 _1964_ (.A(\i_ca.ca_time_const[14] ),
    .B_N(\i_ca.ca_rd_doutb[14] ),
    .X(_0903_));
 sky130_fd_sc_hd__or2b_1 _1965_ (.A(\i_ca.ca_rd_doutb[14] ),
    .B_N(\i_ca.ca_time_const[14] ),
    .X(_0904_));
 sky130_fd_sc_hd__nand2_1 _1966_ (.A(_0903_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__o21bai_1 _1967_ (.A1(\i_ca.ca_time_const[12] ),
    .A2(_0901_),
    .B1_N(_0898_),
    .Y(_0906_));
 sky130_fd_sc_hd__and2b_1 _1968_ (.A_N(_0906_),
    .B(_0895_),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _1969_ (.A(_0899_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__xnor2_1 _1970_ (.A(_0905_),
    .B(_0908_),
    .Y(_0063_));
 sky130_fd_sc_hd__and2b_1 _1971_ (.A_N(\i_ca.ca_rd_doutb[15] ),
    .B(\i_ca.ca_time_const[15] ),
    .X(_0909_));
 sky130_fd_sc_hd__and2b_1 _1972_ (.A_N(\i_ca.ca_time_const[15] ),
    .B(\i_ca.ca_rd_doutb[15] ),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_1 _1973_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__o31a_1 _1974_ (.A1(_0899_),
    .A2(_0905_),
    .A3(_0907_),
    .B1(_0903_),
    .X(_0912_));
 sky130_fd_sc_hd__xnor2_1 _1975_ (.A(_0911_),
    .B(_0912_),
    .Y(_0064_));
 sky130_fd_sc_hd__and3_1 _1976_ (.A(_0903_),
    .B(_0904_),
    .C(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__nand2_1 _1977_ (.A(_0900_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__a211o_1 _1978_ (.A1(_0890_),
    .A2(_0893_),
    .B1(_0914_),
    .C1(_0894_),
    .X(_0915_));
 sky130_fd_sc_hd__and3b_1 _1979_ (.A_N(_0899_),
    .B(_0906_),
    .C(_0913_),
    .X(_0916_));
 sky130_fd_sc_hd__nor2_1 _1980_ (.A(_0910_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__o21a_1 _1981_ (.A1(_0903_),
    .A2(_0909_),
    .B1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__and2_2 _1982_ (.A(_0915_),
    .B(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__xnor2_2 _1983_ (.A(\i_ca.ca_time_const[16] ),
    .B(\i_ca.ca_rd_doutb[16] ),
    .Y(_0920_));
 sky130_fd_sc_hd__xnor2_1 _1984_ (.A(_0919_),
    .B(_0920_),
    .Y(_0065_));
 sky130_fd_sc_hd__and2b_1 _1985_ (.A_N(\i_ca.ca_time_const[17] ),
    .B(\i_ca.ca_rd_doutb[17] ),
    .X(_0921_));
 sky130_fd_sc_hd__and2b_1 _1986_ (.A_N(\i_ca.ca_rd_doutb[17] ),
    .B(\i_ca.ca_time_const[17] ),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_1 _1987_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__or2b_1 _1988_ (.A(\i_ca.ca_time_const[16] ),
    .B_N(\i_ca.ca_rd_doutb[16] ),
    .X(_0924_));
 sky130_fd_sc_hd__or2b_1 _1989_ (.A(_0919_),
    .B_N(_0920_),
    .X(_0925_));
 sky130_fd_sc_hd__and2_1 _1990_ (.A(_0924_),
    .B(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__xnor2_1 _1991_ (.A(_0923_),
    .B(_0926_),
    .Y(_0066_));
 sky130_fd_sc_hd__and2b_1 _1992_ (.A_N(\i_ca.ca_time_const[18] ),
    .B(\i_ca.ca_rd_doutb[18] ),
    .X(_0927_));
 sky130_fd_sc_hd__and2b_1 _1993_ (.A_N(\i_ca.ca_rd_doutb[18] ),
    .B(\i_ca.ca_time_const[18] ),
    .X(_0928_));
 sky130_fd_sc_hd__nor2_1 _1994_ (.A(_0927_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(_0920_),
    .B(_0923_),
    .Y(_0930_));
 sky130_fd_sc_hd__or2_1 _1996_ (.A(_0924_),
    .B(_0922_),
    .X(_0931_));
 sky130_fd_sc_hd__and2b_1 _1997_ (.A_N(_0921_),
    .B(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__o21ai_2 _1998_ (.A1(_0919_),
    .A2(_0930_),
    .B1(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__xor2_1 _1999_ (.A(_0929_),
    .B(_0933_),
    .X(_0067_));
 sky130_fd_sc_hd__xnor2_1 _2000_ (.A(\i_ca.ca_time_const[19] ),
    .B(\i_ca.ca_rd_doutb[19] ),
    .Y(_0934_));
 sky130_fd_sc_hd__a21oi_1 _2001_ (.A1(_0929_),
    .A2(_0933_),
    .B1(_0927_),
    .Y(_0935_));
 sky130_fd_sc_hd__xnor2_1 _2002_ (.A(_0934_),
    .B(_0935_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _2003_ (.A(\i_ca.ca_time_const[19] ),
    .Y(_0936_));
 sky130_fd_sc_hd__o21ai_1 _2004_ (.A1(_0936_),
    .A2(\i_ca.ca_rd_doutb[19] ),
    .B1(\i_ca.ca_rd_doutb[18] ),
    .Y(_0937_));
 sky130_fd_sc_hd__a2bb2o_1 _2005_ (.A1_N(_0937_),
    .A2_N(\i_ca.ca_time_const[18] ),
    .B1(_0936_),
    .B2(\i_ca.ca_rd_doutb[19] ),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_1 _2006_ (.A(_0929_),
    .B(_0934_),
    .Y(_0939_));
 sky130_fd_sc_hd__a211oi_2 _2007_ (.A1(_0915_),
    .A2(_0918_),
    .B1(_0930_),
    .C1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(_0932_),
    .B(_0939_),
    .Y(_0941_));
 sky130_fd_sc_hd__and2b_1 _2009_ (.A_N(\i_ca.ca_time_const[20] ),
    .B(\i_ca.ca_rd_doutb[20] ),
    .X(_0942_));
 sky130_fd_sc_hd__and2b_1 _2010_ (.A_N(\i_ca.ca_rd_doutb[20] ),
    .B(\i_ca.ca_time_const[20] ),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_1 _2011_ (.A(_0942_),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__o31a_1 _2012_ (.A1(_0938_),
    .A2(_0940_),
    .A3(_0941_),
    .B1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__or4_1 _2013_ (.A(_0938_),
    .B(_0940_),
    .C(_0941_),
    .D(_0944_),
    .X(_0946_));
 sky130_fd_sc_hd__and2b_1 _2014_ (.A_N(_0945_),
    .B(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_1 _2015_ (.A(_0947_),
    .X(_0069_));
 sky130_fd_sc_hd__xnor2_1 _2016_ (.A(\i_ca.ca_time_const[21] ),
    .B(\i_ca.ca_rd_doutb[21] ),
    .Y(_0948_));
 sky130_fd_sc_hd__nor2_1 _2017_ (.A(_0942_),
    .B(_0945_),
    .Y(_0949_));
 sky130_fd_sc_hd__xnor2_1 _2018_ (.A(_0948_),
    .B(_0949_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _2019_ (.A(\i_ca.ca_time_const[21] ),
    .Y(_0950_));
 sky130_fd_sc_hd__a21o_1 _2020_ (.A1(_0950_),
    .A2(\i_ca.ca_rd_doutb[21] ),
    .B1(_0942_),
    .X(_0951_));
 sky130_fd_sc_hd__o22a_1 _2021_ (.A1(_0950_),
    .A2(\i_ca.ca_rd_doutb[21] ),
    .B1(_0945_),
    .B2(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__xor2_1 _2022_ (.A(\i_ca.ca_time_const[22] ),
    .B(\i_ca.ca_rd_doutb[22] ),
    .X(_0953_));
 sky130_fd_sc_hd__xnor2_1 _2023_ (.A(_0952_),
    .B(_0953_),
    .Y(_0071_));
 sky130_fd_sc_hd__xor2_1 _2024_ (.A(\i_ca.ca_time_const[0] ),
    .B(\i_ca.ca_time_const[1] ),
    .X(_0049_));
 sky130_fd_sc_hd__and3_1 _2025_ (.A(\i_ca.ca_time_const[0] ),
    .B(\i_ca.ca_time_const[2] ),
    .C(\i_ca.ca_time_const[1] ),
    .X(_0954_));
 sky130_fd_sc_hd__a21oi_1 _2026_ (.A1(\i_ca.ca_time_const[0] ),
    .A2(\i_ca.ca_time_const[1] ),
    .B1(\i_ca.ca_time_const[2] ),
    .Y(_0955_));
 sky130_fd_sc_hd__nor2_1 _2027_ (.A(_0954_),
    .B(_0955_),
    .Y(_0053_));
 sky130_fd_sc_hd__and4_2 _2028_ (.A(\i_ca.ca_time_const[0] ),
    .B(\i_ca.ca_time_const[3] ),
    .C(\i_ca.ca_time_const[2] ),
    .D(\i_ca.ca_time_const[1] ),
    .X(_0956_));
 sky130_fd_sc_hd__nor2_1 _2029_ (.A(\i_ca.ca_time_const[3] ),
    .B(_0954_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_1 _2030_ (.A(_0956_),
    .B(_0957_),
    .Y(_0054_));
 sky130_fd_sc_hd__xor2_1 _2031_ (.A(\i_ca.ca_time_const[4] ),
    .B(_0956_),
    .X(_0055_));
 sky130_fd_sc_hd__and3_2 _2032_ (.A(\i_ca.ca_time_const[5] ),
    .B(\i_ca.ca_time_const[4] ),
    .C(_0956_),
    .X(_0958_));
 sky130_fd_sc_hd__a21oi_1 _2033_ (.A1(\i_ca.ca_time_const[4] ),
    .A2(_0956_),
    .B1(\i_ca.ca_time_const[5] ),
    .Y(_0959_));
 sky130_fd_sc_hd__nor2_1 _2034_ (.A(_0958_),
    .B(_0959_),
    .Y(_0056_));
 sky130_fd_sc_hd__xor2_1 _2035_ (.A(\i_ca.ca_time_const[6] ),
    .B(_0958_),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _2036_ (.A(\i_ca.ca_time_const[7] ),
    .B(\i_ca.ca_time_const[6] ),
    .C(_0958_),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_2 _2037_ (.A(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a21oi_1 _2038_ (.A1(\i_ca.ca_time_const[6] ),
    .A2(_0958_),
    .B1(\i_ca.ca_time_const[7] ),
    .Y(_0962_));
 sky130_fd_sc_hd__nor2_1 _2039_ (.A(_0961_),
    .B(_0962_),
    .Y(_0058_));
 sky130_fd_sc_hd__xor2_1 _2040_ (.A(\i_ca.ca_time_const[8] ),
    .B(_0961_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _2041_ (.A(\i_ca.ca_time_const[9] ),
    .B(\i_ca.ca_time_const[8] ),
    .X(_0963_));
 sky130_fd_sc_hd__nand2_1 _2042_ (.A(_0961_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__a21o_1 _2043_ (.A1(\i_ca.ca_time_const[8] ),
    .A2(_0961_),
    .B1(\i_ca.ca_time_const[9] ),
    .X(_0965_));
 sky130_fd_sc_hd__and2_1 _2044_ (.A(_0964_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_1 _2045_ (.A(_0966_),
    .X(_0060_));
 sky130_fd_sc_hd__xnor2_1 _2046_ (.A(\i_ca.ca_time_const[10] ),
    .B(_0964_),
    .Y(_0039_));
 sky130_fd_sc_hd__a31oi_1 _2047_ (.A1(\i_ca.ca_time_const[10] ),
    .A2(_0961_),
    .A3(_0963_),
    .B1(\i_ca.ca_time_const[11] ),
    .Y(_0967_));
 sky130_fd_sc_hd__and4_2 _2048_ (.A(\i_ca.ca_time_const[11] ),
    .B(\i_ca.ca_time_const[10] ),
    .C(_0961_),
    .D(_0963_),
    .X(_0968_));
 sky130_fd_sc_hd__nor2_1 _2049_ (.A(_0967_),
    .B(_0968_),
    .Y(_0040_));
 sky130_fd_sc_hd__xor2_1 _2050_ (.A(\i_ca.ca_time_const[12] ),
    .B(_0968_),
    .X(_0041_));
 sky130_fd_sc_hd__a21oi_1 _2051_ (.A1(\i_ca.ca_time_const[12] ),
    .A2(_0968_),
    .B1(\i_ca.ca_time_const[13] ),
    .Y(_0969_));
 sky130_fd_sc_hd__and3_2 _2052_ (.A(\i_ca.ca_time_const[13] ),
    .B(\i_ca.ca_time_const[12] ),
    .C(_0968_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_1 _2053_ (.A(_0969_),
    .B(_0970_),
    .Y(_0042_));
 sky130_fd_sc_hd__xor2_1 _2054_ (.A(\i_ca.ca_time_const[14] ),
    .B(_0970_),
    .X(_0043_));
 sky130_fd_sc_hd__a21oi_1 _2055_ (.A1(\i_ca.ca_time_const[14] ),
    .A2(_0970_),
    .B1(\i_ca.ca_time_const[15] ),
    .Y(_0971_));
 sky130_fd_sc_hd__and3_2 _2056_ (.A(\i_ca.ca_time_const[15] ),
    .B(\i_ca.ca_time_const[14] ),
    .C(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_1 _2057_ (.A(_0971_),
    .B(_0972_),
    .Y(_0044_));
 sky130_fd_sc_hd__xor2_1 _2058_ (.A(\i_ca.ca_time_const[16] ),
    .B(_0972_),
    .X(_0045_));
 sky130_fd_sc_hd__a21oi_1 _2059_ (.A1(\i_ca.ca_time_const[16] ),
    .A2(_0972_),
    .B1(\i_ca.ca_time_const[17] ),
    .Y(_0973_));
 sky130_fd_sc_hd__and3_1 _2060_ (.A(\i_ca.ca_time_const[17] ),
    .B(\i_ca.ca_time_const[16] ),
    .C(_0972_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_4 _2061_ (.A(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__nor2_1 _2062_ (.A(_0973_),
    .B(_0975_),
    .Y(_0046_));
 sky130_fd_sc_hd__xor2_1 _2063_ (.A(\i_ca.ca_time_const[18] ),
    .B(_0975_),
    .X(_0047_));
 sky130_fd_sc_hd__a21oi_1 _2064_ (.A1(\i_ca.ca_time_const[18] ),
    .A2(_0975_),
    .B1(\i_ca.ca_time_const[19] ),
    .Y(_0976_));
 sky130_fd_sc_hd__and3_1 _2065_ (.A(\i_ca.ca_time_const[19] ),
    .B(\i_ca.ca_time_const[18] ),
    .C(_0975_),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _2066_ (.A(_0976_),
    .B(_0977_),
    .Y(_0048_));
 sky130_fd_sc_hd__a31o_1 _2067_ (.A1(\i_ca.ca_time_const[19] ),
    .A2(\i_ca.ca_time_const[18] ),
    .A3(_0975_),
    .B1(\i_ca.ca_time_const[20] ),
    .X(_0978_));
 sky130_fd_sc_hd__nand4_4 _2068_ (.A(\i_ca.ca_time_const[19] ),
    .B(\i_ca.ca_time_const[18] ),
    .C(\i_ca.ca_time_const[20] ),
    .D(_0975_),
    .Y(_0979_));
 sky130_fd_sc_hd__and2_1 _2069_ (.A(_0978_),
    .B(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_1 _2070_ (.A(_0980_),
    .X(_0050_));
 sky130_fd_sc_hd__xnor2_1 _2071_ (.A(\i_ca.ca_time_const[21] ),
    .B(_0979_),
    .Y(_0051_));
 sky130_fd_sc_hd__or2_1 _2072_ (.A(_0950_),
    .B(_0979_),
    .X(_0981_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(\i_ca.ca_time_const[22] ),
    .B(_0979_),
    .Y(_0982_));
 sky130_fd_sc_hd__a22o_1 _2074_ (.A1(\i_ca.ca_time_const[22] ),
    .A2(_0981_),
    .B1(_0982_),
    .B2(\i_ca.ca_time_const[21] ),
    .X(_0052_));
 sky130_fd_sc_hd__buf_1 _2075_ (.A(clknet_opt_1_0_wb_clk_i),
    .X(_0983_));
 sky130_fd_sc_hd__buf_1 _2076_ (.A(clknet_1_1__leaf__0983_),
    .X(_0984_));
 sky130_fd_sc_hd__buf_1 _2077_ (.A(clknet_1_1__leaf__0984_),
    .X(_0985_));
 sky130_fd_sc_hd__inv_2 _2079__70 (.A(clknet_1_1__leaf__0985_),
    .Y(net755));
 sky130_fd_sc_hd__inv_2 _2080__71 (.A(clknet_1_1__leaf__0985_),
    .Y(net756));
 sky130_fd_sc_hd__inv_2 _2081__72 (.A(clknet_1_1__leaf__0985_),
    .Y(net757));
 sky130_fd_sc_hd__inv_2 _2082__73 (.A(clknet_1_0__leaf__0985_),
    .Y(net758));
 sky130_fd_sc_hd__inv_2 _2083__74 (.A(clknet_1_1__leaf__0985_),
    .Y(net759));
 sky130_fd_sc_hd__inv_2 _2084__75 (.A(clknet_1_1__leaf__0985_),
    .Y(net760));
 sky130_fd_sc_hd__inv_2 _2085__76 (.A(clknet_1_1__leaf__0985_),
    .Y(net761));
 sky130_fd_sc_hd__inv_2 _2086__77 (.A(clknet_1_0__leaf__0985_),
    .Y(net762));
 sky130_fd_sc_hd__inv_2 _2087__78 (.A(clknet_1_0__leaf__0985_),
    .Y(net763));
 sky130_fd_sc_hd__inv_2 _2089__79 (.A(clknet_1_1__leaf__0986_),
    .Y(net764));
 sky130_fd_sc_hd__buf_1 _2088_ (.A(clknet_1_1__leaf__0984_),
    .X(_0986_));
 sky130_fd_sc_hd__inv_2 _2090__80 (.A(clknet_1_0__leaf__0986_),
    .Y(net765));
 sky130_fd_sc_hd__inv_2 _2091__81 (.A(clknet_1_1__leaf__0986_),
    .Y(net766));
 sky130_fd_sc_hd__inv_2 _2092__82 (.A(clknet_1_0__leaf__0986_),
    .Y(net767));
 sky130_fd_sc_hd__inv_2 _2093__83 (.A(clknet_1_0__leaf__0986_),
    .Y(net768));
 sky130_fd_sc_hd__inv_2 _2094__84 (.A(clknet_1_1__leaf__0986_),
    .Y(net769));
 sky130_fd_sc_hd__inv_2 _2095__85 (.A(clknet_1_0__leaf__0986_),
    .Y(net770));
 sky130_fd_sc_hd__inv_2 _2096__86 (.A(clknet_1_1__leaf__0986_),
    .Y(net771));
 sky130_fd_sc_hd__inv_2 _2097__87 (.A(clknet_1_0__leaf__0986_),
    .Y(net772));
 sky130_fd_sc_hd__inv_2 _2098__88 (.A(clknet_1_1__leaf__0986_),
    .Y(net773));
 sky130_fd_sc_hd__inv_2 _2101__89 (.A(clknet_1_0__leaf__0988_),
    .Y(net774));
 sky130_fd_sc_hd__buf_1 _2099_ (.A(clknet_1_1__leaf__0983_),
    .X(_0987_));
 sky130_fd_sc_hd__buf_1 _2100_ (.A(clknet_1_1_0__0987_),
    .X(_0988_));
 sky130_fd_sc_hd__inv_2 _2102__90 (.A(clknet_1_0__leaf__0988_),
    .Y(net775));
 sky130_fd_sc_hd__inv_2 _2103__91 (.A(clknet_1_1__leaf__0988_),
    .Y(net776));
 sky130_fd_sc_hd__inv_2 _2104__92 (.A(clknet_1_1__leaf__0988_),
    .Y(net777));
 sky130_fd_sc_hd__inv_2 _2105__93 (.A(clknet_1_0__leaf__0988_),
    .Y(net778));
 sky130_fd_sc_hd__inv_2 _2106__94 (.A(clknet_1_1__leaf__0988_),
    .Y(net779));
 sky130_fd_sc_hd__inv_2 _2107__95 (.A(clknet_1_1__leaf__0988_),
    .Y(net780));
 sky130_fd_sc_hd__inv_2 _2108__96 (.A(clknet_1_1__leaf__0988_),
    .Y(net781));
 sky130_fd_sc_hd__inv_2 _2109__97 (.A(clknet_1_0__leaf__0988_),
    .Y(net782));
 sky130_fd_sc_hd__inv_2 _2110__98 (.A(clknet_1_1__leaf__0988_),
    .Y(net783));
 sky130_fd_sc_hd__inv_2 _2112__99 (.A(clknet_1_0__leaf__0989_),
    .Y(net784));
 sky130_fd_sc_hd__buf_1 _2111_ (.A(clknet_1_1_0__0987_),
    .X(_0989_));
 sky130_fd_sc_hd__inv_2 _2113__100 (.A(clknet_1_1__leaf__0989_),
    .Y(net785));
 sky130_fd_sc_hd__inv_2 _2114__101 (.A(clknet_1_0__leaf__0989_),
    .Y(net786));
 sky130_fd_sc_hd__inv_2 _2115__102 (.A(clknet_1_0__leaf__0989_),
    .Y(net787));
 sky130_fd_sc_hd__inv_2 _2116__103 (.A(clknet_1_1__leaf__0989_),
    .Y(net788));
 sky130_fd_sc_hd__inv_2 _2117__104 (.A(clknet_1_1__leaf__0989_),
    .Y(net789));
 sky130_fd_sc_hd__inv_2 _2118__105 (.A(clknet_1_0__leaf__0989_),
    .Y(net790));
 sky130_fd_sc_hd__inv_2 _2119__106 (.A(clknet_1_1__leaf__0989_),
    .Y(net791));
 sky130_fd_sc_hd__inv_2 _2120__107 (.A(clknet_1_0__leaf__0989_),
    .Y(net792));
 sky130_fd_sc_hd__inv_2 _2121__108 (.A(clknet_1_1__leaf__0989_),
    .Y(net793));
 sky130_fd_sc_hd__inv_2 _2123__109 (.A(clknet_1_0__leaf__0990_),
    .Y(net794));
 sky130_fd_sc_hd__buf_1 _2122_ (.A(clknet_1_1_0__0987_),
    .X(_0990_));
 sky130_fd_sc_hd__inv_2 _2124__110 (.A(clknet_1_1__leaf__0990_),
    .Y(net795));
 sky130_fd_sc_hd__inv_2 _2125__111 (.A(clknet_1_0__leaf__0990_),
    .Y(net796));
 sky130_fd_sc_hd__inv_2 _2126__112 (.A(clknet_1_0__leaf__0990_),
    .Y(net797));
 sky130_fd_sc_hd__inv_2 _2127__113 (.A(clknet_1_1__leaf__0990_),
    .Y(net798));
 sky130_fd_sc_hd__inv_2 _2128__114 (.A(clknet_1_1__leaf__0990_),
    .Y(net799));
 sky130_fd_sc_hd__inv_2 _2129__115 (.A(clknet_1_1__leaf__0990_),
    .Y(net800));
 sky130_fd_sc_hd__inv_2 _2130__116 (.A(clknet_1_1__leaf__0990_),
    .Y(net801));
 sky130_fd_sc_hd__inv_2 _2131__117 (.A(clknet_1_0__leaf__0990_),
    .Y(net802));
 sky130_fd_sc_hd__inv_2 _2132__118 (.A(clknet_1_1__leaf__0990_),
    .Y(net803));
 sky130_fd_sc_hd__inv_2 _2134__119 (.A(clknet_1_0__leaf__0991_),
    .Y(net804));
 sky130_fd_sc_hd__buf_1 _2133_ (.A(clknet_1_1_0__0987_),
    .X(_0991_));
 sky130_fd_sc_hd__inv_2 _2135__120 (.A(clknet_1_0__leaf__0991_),
    .Y(net805));
 sky130_fd_sc_hd__inv_2 _2136__121 (.A(clknet_1_0__leaf__0991_),
    .Y(net806));
 sky130_fd_sc_hd__inv_2 _2137__122 (.A(clknet_1_0__leaf__0991_),
    .Y(net807));
 sky130_fd_sc_hd__inv_2 _2138__123 (.A(clknet_1_0__leaf__0991_),
    .Y(net808));
 sky130_fd_sc_hd__inv_2 _2139__124 (.A(clknet_1_1__leaf__0991_),
    .Y(net809));
 sky130_fd_sc_hd__inv_2 _2140__125 (.A(clknet_1_1__leaf__0991_),
    .Y(net810));
 sky130_fd_sc_hd__inv_2 _2141__126 (.A(clknet_1_1__leaf__0991_),
    .Y(net811));
 sky130_fd_sc_hd__inv_2 _2142__127 (.A(clknet_1_1__leaf__0991_),
    .Y(net812));
 sky130_fd_sc_hd__inv_2 _2143__128 (.A(clknet_1_1__leaf__0991_),
    .Y(net813));
 sky130_fd_sc_hd__inv_2 _2145__129 (.A(clknet_1_1__leaf__0992_),
    .Y(net814));
 sky130_fd_sc_hd__buf_1 _2144_ (.A(clknet_1_1_0__0987_),
    .X(_0992_));
 sky130_fd_sc_hd__inv_2 _2146__130 (.A(clknet_1_1__leaf__0992_),
    .Y(net815));
 sky130_fd_sc_hd__inv_2 _2147__131 (.A(clknet_1_0__leaf__0992_),
    .Y(net816));
 sky130_fd_sc_hd__inv_2 _2148__132 (.A(clknet_1_0__leaf__0992_),
    .Y(net817));
 sky130_fd_sc_hd__inv_2 _2149__133 (.A(clknet_1_1__leaf__0992_),
    .Y(net818));
 sky130_fd_sc_hd__inv_2 _2150__134 (.A(clknet_1_1__leaf__0992_),
    .Y(net819));
 sky130_fd_sc_hd__inv_2 _2151__135 (.A(clknet_1_1__leaf__0992_),
    .Y(net820));
 sky130_fd_sc_hd__inv_2 _2152__136 (.A(clknet_1_0__leaf__0992_),
    .Y(net821));
 sky130_fd_sc_hd__inv_2 _2153__137 (.A(clknet_1_0__leaf__0992_),
    .Y(net822));
 sky130_fd_sc_hd__inv_2 _2154__138 (.A(clknet_1_0__leaf__0992_),
    .Y(net823));
 sky130_fd_sc_hd__inv_2 _2156__139 (.A(clknet_1_1__leaf__0993_),
    .Y(net824));
 sky130_fd_sc_hd__buf_1 _2155_ (.A(clknet_1_1_0__0987_),
    .X(_0993_));
 sky130_fd_sc_hd__inv_2 _2157__140 (.A(clknet_1_0__leaf__0993_),
    .Y(net825));
 sky130_fd_sc_hd__inv_2 _2158__141 (.A(clknet_1_1__leaf__0993_),
    .Y(net826));
 sky130_fd_sc_hd__inv_2 _2159__142 (.A(clknet_1_0__leaf__0993_),
    .Y(net827));
 sky130_fd_sc_hd__inv_2 _2160__143 (.A(clknet_1_0__leaf__0993_),
    .Y(net828));
 sky130_fd_sc_hd__inv_2 _2161__144 (.A(clknet_1_0__leaf__0993_),
    .Y(net829));
 sky130_fd_sc_hd__inv_2 _2162__145 (.A(clknet_1_1__leaf__0993_),
    .Y(net830));
 sky130_fd_sc_hd__inv_2 _2163__146 (.A(clknet_1_1__leaf__0993_),
    .Y(net831));
 sky130_fd_sc_hd__inv_2 _2164__147 (.A(clknet_1_1__leaf__0993_),
    .Y(net832));
 sky130_fd_sc_hd__inv_2 _2165__148 (.A(clknet_1_1__leaf__0993_),
    .Y(net833));
 sky130_fd_sc_hd__inv_2 _2167__149 (.A(clknet_1_1__leaf__0994_),
    .Y(net834));
 sky130_fd_sc_hd__buf_1 _2166_ (.A(clknet_1_0_0__0987_),
    .X(_0994_));
 sky130_fd_sc_hd__inv_2 _2217__150 (.A(clknet_1_1__leaf__0994_),
    .Y(net835));
 sky130_fd_sc_hd__nand2b_4 _2168_ (.A_N(net331),
    .B(\i_ca.hs_ready_meta ),
    .Y(_0995_));
 sky130_fd_sc_hd__clkbuf_8 _2169_ (.A(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _2170_ (.A0(\i_ca.ca_time_const[0] ),
    .A1(net308),
    .S(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _2171_ (.A(_0997_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2172_ (.A0(\i_ca.ca_time_const[1] ),
    .A1(net319),
    .S(_0996_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _2173_ (.A(_0998_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(\i_ca.ca_time_const[2] ),
    .A1(net323),
    .S(_0996_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_1 _2175_ (.A(_0999_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(\i_ca.ca_time_const[3] ),
    .A1(net324),
    .S(_0996_),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_1 _2177_ (.A(_1000_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2178_ (.A0(\i_ca.ca_time_const[4] ),
    .A1(net325),
    .S(_0996_),
    .X(_1001_));
 sky130_fd_sc_hd__clkbuf_1 _2179_ (.A(_1001_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2180_ (.A0(\i_ca.ca_time_const[5] ),
    .A1(net326),
    .S(_0996_),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_1 _2181_ (.A(_1002_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(\i_ca.ca_time_const[6] ),
    .A1(net327),
    .S(_0996_),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_1 _2183_ (.A(_1003_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2184_ (.A0(\i_ca.ca_time_const[7] ),
    .A1(net328),
    .S(_0996_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_1 _2185_ (.A(_1004_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2186_ (.A0(\i_ca.ca_time_const[8] ),
    .A1(net329),
    .S(_0996_),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _2187_ (.A(_1005_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(\i_ca.ca_time_const[9] ),
    .A1(net330),
    .S(_0996_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _2189_ (.A(_1006_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_8 _2190_ (.A(_0995_),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _2191_ (.A0(\i_ca.ca_time_const[10] ),
    .A1(net309),
    .S(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_1 _2192_ (.A(_1008_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2193_ (.A0(\i_ca.ca_time_const[11] ),
    .A1(net310),
    .S(_1007_),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _2194_ (.A(_1009_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _2195_ (.A0(\i_ca.ca_time_const[12] ),
    .A1(net311),
    .S(_1007_),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _2196_ (.A(_1010_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(\i_ca.ca_time_const[13] ),
    .A1(net312),
    .S(_1007_),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _2198_ (.A(_1011_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(\i_ca.ca_time_const[14] ),
    .A1(net313),
    .S(_1007_),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _2200_ (.A(_1012_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(\i_ca.ca_time_const[15] ),
    .A1(net314),
    .S(_1007_),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _2202_ (.A(_1013_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(\i_ca.ca_time_const[16] ),
    .A1(net315),
    .S(_1007_),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _2204_ (.A(_1014_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _2205_ (.A0(\i_ca.ca_time_const[17] ),
    .A1(net316),
    .S(_1007_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _2206_ (.A(_1015_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(\i_ca.ca_time_const[18] ),
    .A1(net317),
    .S(_1007_),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _2208_ (.A(_1016_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(\i_ca.ca_time_const[19] ),
    .A1(net318),
    .S(_1007_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _2210_ (.A(_1017_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(\i_ca.ca_time_const[20] ),
    .A1(net320),
    .S(_0995_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _2212_ (.A(_1018_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(\i_ca.ca_time_const[21] ),
    .A1(net321),
    .S(_0995_),
    .X(_1019_));
 sky130_fd_sc_hd__clkbuf_1 _2214_ (.A(_1019_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(\i_ca.ca_time_const[22] ),
    .A1(net322),
    .S(_0995_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _2216_ (.A(_1020_),
    .X(_0374_));
 sky130_fd_sc_hd__inv_2 _2218__151 (.A(clknet_1_1__leaf__0994_),
    .Y(net836));
 sky130_fd_sc_hd__inv_2 _2219__152 (.A(clknet_1_1__leaf__0994_),
    .Y(net837));
 sky130_fd_sc_hd__inv_2 _2220__153 (.A(clknet_1_0__leaf__0994_),
    .Y(net838));
 sky130_fd_sc_hd__inv_2 _2221__154 (.A(clknet_1_0__leaf__0994_),
    .Y(net839));
 sky130_fd_sc_hd__inv_2 _2222__155 (.A(clknet_1_0__leaf__0994_),
    .Y(net840));
 sky130_fd_sc_hd__inv_2 _2223__156 (.A(clknet_1_0__leaf__0994_),
    .Y(net841));
 sky130_fd_sc_hd__inv_2 _2224__157 (.A(clknet_1_0__leaf__0994_),
    .Y(net842));
 sky130_fd_sc_hd__inv_2 _2225__158 (.A(clknet_1_0__leaf__0994_),
    .Y(net843));
 sky130_fd_sc_hd__inv_2 _2227__159 (.A(clknet_1_1__leaf__1021_),
    .Y(net844));
 sky130_fd_sc_hd__buf_1 _2226_ (.A(clknet_1_0_0__0987_),
    .X(_1021_));
 sky130_fd_sc_hd__inv_2 _2228__160 (.A(clknet_1_1__leaf__1021_),
    .Y(net845));
 sky130_fd_sc_hd__inv_2 _2229__161 (.A(clknet_1_0__leaf__1021_),
    .Y(net846));
 sky130_fd_sc_hd__inv_2 _2230__162 (.A(clknet_1_0__leaf__1021_),
    .Y(net847));
 sky130_fd_sc_hd__inv_2 _2231__163 (.A(clknet_1_0__leaf__1021_),
    .Y(net848));
 sky130_fd_sc_hd__inv_2 _2232__164 (.A(clknet_1_0__leaf__1021_),
    .Y(net849));
 sky130_fd_sc_hd__inv_2 _2233__165 (.A(clknet_1_0__leaf__1021_),
    .Y(net850));
 sky130_fd_sc_hd__inv_2 _2234__166 (.A(clknet_1_1__leaf__1021_),
    .Y(net851));
 sky130_fd_sc_hd__inv_2 _2235__167 (.A(clknet_1_1__leaf__1021_),
    .Y(net852));
 sky130_fd_sc_hd__inv_2 _2236__168 (.A(clknet_1_1__leaf__1021_),
    .Y(net853));
 sky130_fd_sc_hd__inv_2 _2238__169 (.A(clknet_1_0__leaf__1022_),
    .Y(net854));
 sky130_fd_sc_hd__buf_1 _2237_ (.A(clknet_1_0_0__0987_),
    .X(_1022_));
 sky130_fd_sc_hd__inv_2 _2239__170 (.A(clknet_1_0__leaf__1022_),
    .Y(net855));
 sky130_fd_sc_hd__inv_2 _2240__171 (.A(clknet_1_0__leaf__1022_),
    .Y(net856));
 sky130_fd_sc_hd__inv_2 _2241__172 (.A(clknet_1_0__leaf__1022_),
    .Y(net857));
 sky130_fd_sc_hd__inv_2 _2242__173 (.A(clknet_1_0__leaf__1022_),
    .Y(net858));
 sky130_fd_sc_hd__inv_2 _2243__174 (.A(clknet_1_1__leaf__1022_),
    .Y(net859));
 sky130_fd_sc_hd__inv_2 _2244__175 (.A(clknet_1_1__leaf__1022_),
    .Y(net860));
 sky130_fd_sc_hd__inv_2 _2245__176 (.A(clknet_1_1__leaf__1022_),
    .Y(net861));
 sky130_fd_sc_hd__inv_2 _2246__177 (.A(clknet_1_1__leaf__1022_),
    .Y(net862));
 sky130_fd_sc_hd__inv_2 _2247__178 (.A(clknet_1_1__leaf__1022_),
    .Y(net863));
 sky130_fd_sc_hd__inv_2 _2249__179 (.A(clknet_1_0__leaf__1023_),
    .Y(net864));
 sky130_fd_sc_hd__buf_1 _2248_ (.A(clknet_1_0_0__0987_),
    .X(_1023_));
 sky130_fd_sc_hd__inv_2 _2250__180 (.A(clknet_1_0__leaf__1023_),
    .Y(net865));
 sky130_fd_sc_hd__inv_2 _2251__181 (.A(clknet_1_0__leaf__1023_),
    .Y(net866));
 sky130_fd_sc_hd__inv_2 _2252__182 (.A(clknet_1_0__leaf__1023_),
    .Y(net867));
 sky130_fd_sc_hd__inv_2 _2253__183 (.A(clknet_1_0__leaf__1023_),
    .Y(net868));
 sky130_fd_sc_hd__inv_2 _2254__184 (.A(clknet_1_1__leaf__1023_),
    .Y(net869));
 sky130_fd_sc_hd__inv_2 _2255__185 (.A(clknet_1_1__leaf__1023_),
    .Y(net870));
 sky130_fd_sc_hd__inv_2 _2256__186 (.A(clknet_1_1__leaf__1023_),
    .Y(net871));
 sky130_fd_sc_hd__inv_2 _2257__187 (.A(clknet_1_1__leaf__1023_),
    .Y(net872));
 sky130_fd_sc_hd__inv_2 _2258__188 (.A(clknet_1_1__leaf__1023_),
    .Y(net873));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__buf_1 _2259_ (.A(clknet_1_0__leaf__0983_),
    .X(_1024_));
 sky130_fd_sc_hd__inv_2 _2261__10 (.A(clknet_1_1__leaf__1024_),
    .Y(net695));
 sky130_fd_sc_hd__inv_2 _2262__11 (.A(clknet_1_1__leaf__1024_),
    .Y(net696));
 sky130_fd_sc_hd__inv_2 _2263__12 (.A(clknet_1_1__leaf__1024_),
    .Y(net697));
 sky130_fd_sc_hd__inv_2 _2264__13 (.A(clknet_1_0__leaf__1024_),
    .Y(net698));
 sky130_fd_sc_hd__inv_2 _2265__14 (.A(clknet_1_0__leaf__1024_),
    .Y(net699));
 sky130_fd_sc_hd__inv_2 _2266__15 (.A(clknet_1_0__leaf__1024_),
    .Y(net700));
 sky130_fd_sc_hd__inv_2 _2267__16 (.A(clknet_1_0__leaf__1024_),
    .Y(net701));
 sky130_fd_sc_hd__inv_2 _2268__17 (.A(clknet_1_0__leaf__1024_),
    .Y(net702));
 sky130_fd_sc_hd__inv_2 _2269__18 (.A(clknet_1_1__leaf__1024_),
    .Y(net703));
 sky130_fd_sc_hd__inv_2 _2271__19 (.A(clknet_1_0__leaf__1025_),
    .Y(net704));
 sky130_fd_sc_hd__buf_1 _2270_ (.A(clknet_1_0__leaf__0983_),
    .X(_1025_));
 sky130_fd_sc_hd__inv_2 _2272__20 (.A(clknet_1_1__leaf__1025_),
    .Y(net705));
 sky130_fd_sc_hd__inv_2 _2273__21 (.A(clknet_1_0__leaf__1025_),
    .Y(net706));
 sky130_fd_sc_hd__inv_2 _2274__22 (.A(clknet_1_0__leaf__1025_),
    .Y(net707));
 sky130_fd_sc_hd__inv_2 _2275__23 (.A(clknet_1_1__leaf__1025_),
    .Y(net708));
 sky130_fd_sc_hd__inv_2 _2276__24 (.A(clknet_1_1__leaf__1025_),
    .Y(net709));
 sky130_fd_sc_hd__inv_2 _2277__25 (.A(clknet_1_1__leaf__1025_),
    .Y(net710));
 sky130_fd_sc_hd__inv_2 _2278__26 (.A(clknet_1_0__leaf__1025_),
    .Y(net711));
 sky130_fd_sc_hd__inv_2 _2279__27 (.A(clknet_1_1__leaf__1025_),
    .Y(net712));
 sky130_fd_sc_hd__inv_2 _2280__28 (.A(clknet_1_0__leaf__1025_),
    .Y(net713));
 sky130_fd_sc_hd__inv_2 _2282__29 (.A(clknet_1_1__leaf__1026_),
    .Y(net714));
 sky130_fd_sc_hd__buf_1 _2281_ (.A(clknet_1_0__leaf__0983_),
    .X(_1026_));
 sky130_fd_sc_hd__inv_2 _2283__30 (.A(clknet_1_0__leaf__1026_),
    .Y(net715));
 sky130_fd_sc_hd__inv_2 _2284__31 (.A(clknet_1_1__leaf__1026_),
    .Y(net716));
 sky130_fd_sc_hd__inv_2 _2285__32 (.A(clknet_1_1__leaf__1026_),
    .Y(net717));
 sky130_fd_sc_hd__inv_2 _2286__33 (.A(clknet_1_0__leaf__1026_),
    .Y(net718));
 sky130_fd_sc_hd__inv_2 _2287__34 (.A(clknet_1_0__leaf__1026_),
    .Y(net719));
 sky130_fd_sc_hd__inv_2 _2288__35 (.A(clknet_1_0__leaf__1026_),
    .Y(net720));
 sky130_fd_sc_hd__inv_2 _2289__36 (.A(clknet_1_0__leaf__1026_),
    .Y(net721));
 sky130_fd_sc_hd__inv_2 _2290__37 (.A(clknet_1_1__leaf__1026_),
    .Y(net722));
 sky130_fd_sc_hd__inv_2 _2291__38 (.A(clknet_1_1__leaf__1026_),
    .Y(net723));
 sky130_fd_sc_hd__inv_2 _2293__39 (.A(clknet_1_1__leaf__1027_),
    .Y(net724));
 sky130_fd_sc_hd__buf_1 _2292_ (.A(clknet_1_0__leaf__0983_),
    .X(_1027_));
 sky130_fd_sc_hd__inv_2 _2294__40 (.A(clknet_1_1__leaf__1027_),
    .Y(net725));
 sky130_fd_sc_hd__inv_2 _2295__41 (.A(clknet_1_0__leaf__1027_),
    .Y(net726));
 sky130_fd_sc_hd__inv_2 _2296__42 (.A(clknet_1_0__leaf__1027_),
    .Y(net727));
 sky130_fd_sc_hd__inv_2 _2297__43 (.A(clknet_1_0__leaf__1027_),
    .Y(net728));
 sky130_fd_sc_hd__inv_2 _2298__44 (.A(clknet_1_0__leaf__1027_),
    .Y(net729));
 sky130_fd_sc_hd__inv_2 _2299__45 (.A(clknet_1_0__leaf__1027_),
    .Y(net730));
 sky130_fd_sc_hd__inv_2 _2300__46 (.A(clknet_1_0__leaf__1027_),
    .Y(net731));
 sky130_fd_sc_hd__inv_2 _2301__47 (.A(clknet_1_1__leaf__1027_),
    .Y(net732));
 sky130_fd_sc_hd__inv_2 _2302__48 (.A(clknet_1_1__leaf__1027_),
    .Y(net733));
 sky130_fd_sc_hd__inv_2 _2304__49 (.A(clknet_1_1__leaf__1028_),
    .Y(net734));
 sky130_fd_sc_hd__buf_1 _2303_ (.A(clknet_1_1__leaf__0983_),
    .X(_1028_));
 sky130_fd_sc_hd__inv_2 _2305__50 (.A(clknet_1_1__leaf__1028_),
    .Y(net735));
 sky130_fd_sc_hd__inv_2 _2306__51 (.A(clknet_1_0__leaf__1028_),
    .Y(net736));
 sky130_fd_sc_hd__inv_2 _2307__52 (.A(clknet_1_0__leaf__1028_),
    .Y(net737));
 sky130_fd_sc_hd__inv_2 _2308__53 (.A(clknet_1_0__leaf__1028_),
    .Y(net738));
 sky130_fd_sc_hd__inv_2 _2309__54 (.A(clknet_1_0__leaf__1028_),
    .Y(net739));
 sky130_fd_sc_hd__inv_2 _2310__55 (.A(clknet_1_1__leaf__1028_),
    .Y(net740));
 sky130_fd_sc_hd__inv_2 _2311__56 (.A(clknet_1_1__leaf__1028_),
    .Y(net741));
 sky130_fd_sc_hd__inv_2 _2312__57 (.A(clknet_1_1__leaf__1028_),
    .Y(net742));
 sky130_fd_sc_hd__inv_2 _2313__58 (.A(clknet_1_0__leaf__1028_),
    .Y(net743));
 sky130_fd_sc_hd__inv_2 _2315__59 (.A(clknet_1_0__leaf__1029_),
    .Y(net744));
 sky130_fd_sc_hd__buf_1 _2314_ (.A(clknet_1_1__leaf__0983_),
    .X(_1029_));
 sky130_fd_sc_hd__inv_2 _2316__60 (.A(clknet_1_0__leaf__1029_),
    .Y(net745));
 sky130_fd_sc_hd__inv_2 _2317__61 (.A(clknet_1_0__leaf__1029_),
    .Y(net746));
 sky130_fd_sc_hd__inv_2 _2318__62 (.A(clknet_1_1__leaf__1029_),
    .Y(net747));
 sky130_fd_sc_hd__inv_2 _2319__63 (.A(clknet_1_0__leaf__1029_),
    .Y(net748));
 sky130_fd_sc_hd__inv_2 _2320__64 (.A(clknet_1_1__leaf__1029_),
    .Y(net749));
 sky130_fd_sc_hd__inv_2 _2321__65 (.A(clknet_1_0__leaf__1029_),
    .Y(net750));
 sky130_fd_sc_hd__inv_2 _2322__66 (.A(clknet_1_1__leaf__1029_),
    .Y(net751));
 sky130_fd_sc_hd__inv_2 _2323__67 (.A(clknet_1_1__leaf__1029_),
    .Y(net752));
 sky130_fd_sc_hd__inv_2 _2324__68 (.A(clknet_1_1__leaf__1029_),
    .Y(net753));
 sky130_fd_sc_hd__inv_2 _2078__69 (.A(clknet_1_0__leaf__0985_),
    .Y(net754));
 sky130_fd_sc_hd__inv_2 _2326__2 (.A(clknet_1_0__leaf__0984_),
    .Y(net687));
 sky130_fd_sc_hd__inv_2 _2327__3 (.A(clknet_1_0__leaf__0984_),
    .Y(net688));
 sky130_fd_sc_hd__inv_2 _2328__4 (.A(clknet_1_0__leaf__0984_),
    .Y(net689));
 sky130_fd_sc_hd__inv_2 _2329__5 (.A(clknet_1_0__leaf__0984_),
    .Y(net690));
 sky130_fd_sc_hd__inv_2 _2330__6 (.A(clknet_1_0__leaf__0984_),
    .Y(net691));
 sky130_fd_sc_hd__inv_2 _2331__7 (.A(clknet_1_0__leaf__0984_),
    .Y(net692));
 sky130_fd_sc_hd__inv_2 _2332__8 (.A(clknet_1_1__leaf__0984_),
    .Y(net693));
 sky130_fd_sc_hd__inv_2 _2260__9 (.A(clknet_1_0__leaf__1024_),
    .Y(net694));
 sky130_fd_sc_hd__inv_2 _2333_ (.A(_0761_),
    .Y(_1030_));
 sky130_fd_sc_hd__and2_1 _2334_ (.A(_1030_),
    .B(_0858_),
    .X(_1031_));
 sky130_fd_sc_hd__or2_1 _2335_ (.A(\i_ca.ca_wr_fsm_state[7] ),
    .B(\i_ca.ca_wr_fsm_state[16] ),
    .X(_1032_));
 sky130_fd_sc_hd__buf_4 _2336_ (.A(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__or2_4 _2337_ (.A(\i_ca.ca_wr_fsm_state[4] ),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__nor2_1 _2338_ (.A(\i_ca.ca_wr_fsm_state[1] ),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__nand2_1 _2339_ (.A(_0764_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__and4b_2 _2340_ (.A_N(_0721_),
    .B(_0842_),
    .C(_1031_),
    .D(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__and2_1 _2341_ (.A(\i_ca.ca_wr_add_fill[1] ),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__or2_1 _2342_ (.A(\i_ca.ca_wr_fsm_state[1] ),
    .B(_1034_),
    .X(_1039_));
 sky130_fd_sc_hd__a21oi_1 _2343_ (.A1(_1039_),
    .A2(_1037_),
    .B1(\i_ca.ca_wr_add_fill[1] ),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_1 _2344_ (.A(_1038_),
    .B(_1040_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_2 _2345_ (.A(_1035_),
    .B(_1037_),
    .Y(_1041_));
 sky130_fd_sc_hd__and3_1 _2346_ (.A(\i_ca.ca_wr_add_fill[1] ),
    .B(\i_ca.ca_wr_add_fill[2] ),
    .C(_1037_),
    .X(_1042_));
 sky130_fd_sc_hd__inv_2 _2347_ (.A(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__o211a_1 _2348_ (.A1(\i_ca.ca_wr_add_fill[2] ),
    .A2(_1038_),
    .B1(_1041_),
    .C1(_1043_),
    .X(_0418_));
 sky130_fd_sc_hd__and4_2 _2349_ (.A(\i_ca.ca_wr_add_fill[1] ),
    .B(\i_ca.ca_wr_add_fill[3] ),
    .C(\i_ca.ca_wr_add_fill[2] ),
    .D(_1037_),
    .X(_1044_));
 sky130_fd_sc_hd__inv_2 _2350_ (.A(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__o211a_1 _2351_ (.A1(\i_ca.ca_wr_add_fill[3] ),
    .A2(_1042_),
    .B1(_1045_),
    .C1(_1041_),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _2352_ (.A(\i_ca.ca_wr_add_fill[4] ),
    .B(_1044_),
    .X(_1046_));
 sky130_fd_sc_hd__nor2_1 _2353_ (.A(\i_ca.ca_wr_add_fill[4] ),
    .B(_1044_),
    .Y(_1047_));
 sky130_fd_sc_hd__or4bb_1 _2354_ (.A(\i_ca.ca_wr_add_fill[8] ),
    .B(\i_ca.ca_wr_add_fill[6] ),
    .C_N(\i_ca.ca_wr_add_fill[4] ),
    .D_N(\i_ca.ca_wr_add_fill[5] ),
    .X(_1048_));
 sky130_fd_sc_hd__o21ai_1 _2355_ (.A1(\i_ca.ca_wr_add_fill[7] ),
    .A2(_1048_),
    .B1(_1039_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand2_1 _2356_ (.A(_1037_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__o21ai_1 _2357_ (.A1(_1046_),
    .A2(_1047_),
    .B1(_1050_),
    .Y(_0420_));
 sky130_fd_sc_hd__and3_1 _2358_ (.A(\i_ca.ca_wr_add_fill[5] ),
    .B(\i_ca.ca_wr_add_fill[4] ),
    .C(_1044_),
    .X(_1051_));
 sky130_fd_sc_hd__o21ai_1 _2359_ (.A1(\i_ca.ca_wr_add_fill[5] ),
    .A2(_1046_),
    .B1(_1041_),
    .Y(_1052_));
 sky130_fd_sc_hd__nor2_1 _2360_ (.A(_1051_),
    .B(_1052_),
    .Y(_0421_));
 sky130_fd_sc_hd__and2_1 _2361_ (.A(\i_ca.ca_wr_add_fill[6] ),
    .B(_1051_),
    .X(_1053_));
 sky130_fd_sc_hd__inv_2 _2362_ (.A(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__o211a_1 _2363_ (.A1(\i_ca.ca_wr_add_fill[6] ),
    .A2(_1051_),
    .B1(_1054_),
    .C1(_1050_),
    .X(_0422_));
 sky130_fd_sc_hd__a21boi_1 _2364_ (.A1(\i_ca.ca_wr_add_fill[7] ),
    .A2(_1053_),
    .B1_N(_1041_),
    .Y(_1055_));
 sky130_fd_sc_hd__o21a_1 _2365_ (.A1(\i_ca.ca_wr_add_fill[7] ),
    .A2(_1053_),
    .B1(_1055_),
    .X(_0423_));
 sky130_fd_sc_hd__nor2_1 _2366_ (.A(\i_ca.ca_wr_add_fill[8] ),
    .B(_1035_),
    .Y(_1056_));
 sky130_fd_sc_hd__a31o_1 _2367_ (.A1(\i_ca.ca_wr_add_fill[7] ),
    .A2(\i_ca.ca_wr_add_fill[6] ),
    .A3(_1051_),
    .B1(\i_ca.ca_wr_add_fill[8] ),
    .X(_1057_));
 sky130_fd_sc_hd__o21a_1 _2368_ (.A1(_1055_),
    .A2(_1056_),
    .B1(_1057_),
    .X(_0424_));
 sky130_fd_sc_hd__and2_1 _2369_ (.A(_0720_),
    .B(\i_ca.ca_rd_doutb[23] ),
    .X(_1058_));
 sky130_fd_sc_hd__or2_4 _2370_ (.A(_0719_),
    .B(_1033_),
    .X(_1059_));
 sky130_fd_sc_hd__buf_4 _2371_ (.A(\i_ca.ca_wr_fsm_state[7] ),
    .X(_1060_));
 sky130_fd_sc_hd__nor2_1 _2372_ (.A(_1060_),
    .B(\i_ca.ca_wr_fsm_state[16] ),
    .Y(_1061_));
 sky130_fd_sc_hd__or2_2 _2373_ (.A(\i_ca.ca_wr_com_const ),
    .B(_0704_),
    .X(_1062_));
 sky130_fd_sc_hd__nor2_1 _2374_ (.A(_0718_),
    .B(\i_ca.ca_rd_doutb_31_23 ),
    .Y(_1063_));
 sky130_fd_sc_hd__o21ai_1 _2375_ (.A1(_1062_),
    .A2(_1063_),
    .B1(_0719_),
    .Y(_1064_));
 sky130_fd_sc_hd__or2_1 _2376_ (.A(\i_ca.ca_wr_sync_update ),
    .B(_0706_),
    .X(_1065_));
 sky130_fd_sc_hd__o2111a_1 _2377_ (.A1(_0708_),
    .A2(_1061_),
    .B1(_1064_),
    .C1(_1065_),
    .D1(_1030_),
    .X(_1066_));
 sky130_fd_sc_hd__o211ai_4 _2378_ (.A1(\i_ca.ca_wr_fsm_state[0] ),
    .A2(_1059_),
    .B1(_1066_),
    .C1(_0858_),
    .Y(_1067_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(_1058_),
    .A1(\i_ca.ca_wr_add_start[0] ),
    .S(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _2380_ (.A(_1068_),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _2381_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[24] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[1] ),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_4 _2382_ (.A(\i_ca.ca_wr_add_start[1] ),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(_1069_),
    .A1(_1070_),
    .S(_1067_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_1071_),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _2385_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[25] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[2] ),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _2386_ (.A0(_1072_),
    .A1(\i_ca.ca_wr_add_start[2] ),
    .S(_1067_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _2387_ (.A(_1073_),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _2388_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[26] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[3] ),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(_1074_),
    .A1(\i_ca.ca_wr_add_start[3] ),
    .S(_1067_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_1075_),
    .X(_0428_));
 sky130_fd_sc_hd__a21bo_1 _2391_ (.A1(\i_ca.ca_wr_add_fill[4] ),
    .A2(_1033_),
    .B1_N(_1059_),
    .X(_1076_));
 sky130_fd_sc_hd__a21o_1 _2392_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[27] ),
    .B1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(_1077_),
    .A1(\i_ca.ca_wr_add_start[4] ),
    .S(_1067_),
    .X(_1078_));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(_1078_),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _2395_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[28] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[5] ),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(_1079_),
    .A1(\i_ca.ca_wr_add_start[5] ),
    .S(_1067_),
    .X(_1080_));
 sky130_fd_sc_hd__clkbuf_1 _2397_ (.A(_1080_),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _2398_ (.A1(_0720_),
    .A2(\i_ca.ca_rd_doutb[29] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[6] ),
    .X(_1081_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(_1081_),
    .A1(\i_ca.ca_wr_add_start[6] ),
    .S(_1067_),
    .X(_1082_));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(_1082_),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _2401_ (.A1(_0719_),
    .A2(\i_ca.ca_rd_doutb[30] ),
    .B1(_1033_),
    .B2(\i_ca.ca_wr_add_fill[7] ),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(_1083_),
    .A1(\i_ca.ca_wr_add_start[7] ),
    .S(_1067_),
    .X(_1084_));
 sky130_fd_sc_hd__clkbuf_1 _2403_ (.A(_1084_),
    .X(_0432_));
 sky130_fd_sc_hd__buf_4 _2404_ (.A(_1061_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_1 _2405_ (.A(_1085_),
    .B(_1067_),
    .Y(_1086_));
 sky130_fd_sc_hd__a22o_1 _2406_ (.A1(\i_ca.ca_wr_add_start[8] ),
    .A2(_1067_),
    .B1(_1086_),
    .B2(\i_ca.ca_wr_add_fill[8] ),
    .X(_0433_));
 sky130_fd_sc_hd__nor3_4 _2407_ (.A(\i_ca.ca_wr_fsm_state[3] ),
    .B(\i_ca.ca_wr_fsm_state[15] ),
    .C(_1034_),
    .Y(_1087_));
 sky130_fd_sc_hd__buf_4 _2408_ (.A(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__or3_4 _2409_ (.A(\i_ca.ca_wr_fsm_state[16] ),
    .B(\i_ca.ca_wr_fsm_state[4] ),
    .C(_0711_),
    .X(_1089_));
 sky130_fd_sc_hd__buf_4 _2410_ (.A(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__or3_4 _2411_ (.A(\i_ca.ca_wr_fsm_state[3] ),
    .B(\i_ca.ca_wr_fsm_state[15] ),
    .C(_0001_),
    .X(_1091_));
 sky130_fd_sc_hd__clkbuf_4 _2412_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__and2_1 _2413_ (.A(\i_ca.ca_wr_douta[0] ),
    .B(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__a221o_1 _2414_ (.A1(\i_ca.hs_write_dbus_wr_data_const[0] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[0] ),
    .C1(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__o41a_2 _2415_ (.A1(_0719_),
    .A2(\i_ca.ca_wr_fsm_state[3] ),
    .A3(\i_ca.ca_wr_fsm_state[15] ),
    .A4(_1034_),
    .B1(_0842_),
    .X(_1095_));
 sky130_fd_sc_hd__and3_4 _2416_ (.A(_0705_),
    .B(_0858_),
    .C(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__buf_4 _2417_ (.A(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(\i_ca.ca_wr_dina[0] ),
    .A1(_1094_),
    .S(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__clkbuf_1 _2419_ (.A(_1098_),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _2420_ (.A(\i_ca.ca_wr_douta[1] ),
    .B(_1092_),
    .X(_1099_));
 sky130_fd_sc_hd__a221o_1 _2421_ (.A1(\i_ca.hs_write_dbus_wr_data_const[1] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[1] ),
    .C1(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(\i_ca.ca_wr_dina[1] ),
    .A1(_1100_),
    .S(_1097_),
    .X(_1101_));
 sky130_fd_sc_hd__clkbuf_1 _2423_ (.A(_1101_),
    .X(_0435_));
 sky130_fd_sc_hd__and2_1 _2424_ (.A(\i_ca.ca_wr_douta[2] ),
    .B(_1092_),
    .X(_1102_));
 sky130_fd_sc_hd__a221o_1 _2425_ (.A1(\i_ca.hs_write_dbus_wr_data_const[2] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[2] ),
    .C1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(\i_ca.ca_wr_dina[2] ),
    .A1(_1103_),
    .S(_1097_),
    .X(_1104_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_1104_),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _2428_ (.A(\i_ca.ca_wr_douta[3] ),
    .B(_1092_),
    .X(_1105_));
 sky130_fd_sc_hd__a221o_1 _2429_ (.A1(\i_ca.hs_write_dbus_wr_data_const[3] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[3] ),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(\i_ca.ca_wr_dina[3] ),
    .A1(_1106_),
    .S(_1097_),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _2431_ (.A(_1107_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _2432_ (.A(\i_ca.ca_wr_douta[4] ),
    .B(_1092_),
    .X(_1108_));
 sky130_fd_sc_hd__a221o_1 _2433_ (.A1(\i_ca.hs_write_dbus_wr_data_const[4] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[4] ),
    .C1(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(\i_ca.ca_wr_dina[4] ),
    .A1(_1109_),
    .S(_1097_),
    .X(_1110_));
 sky130_fd_sc_hd__clkbuf_1 _2435_ (.A(_1110_),
    .X(_0438_));
 sky130_fd_sc_hd__and2_1 _2436_ (.A(\i_ca.ca_wr_douta[5] ),
    .B(_1092_),
    .X(_1111_));
 sky130_fd_sc_hd__a221o_1 _2437_ (.A1(\i_ca.hs_write_dbus_wr_data_const[5] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[5] ),
    .C1(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\i_ca.ca_wr_dina[5] ),
    .A1(_1112_),
    .S(_1097_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_1113_),
    .X(_0439_));
 sky130_fd_sc_hd__and2_1 _2440_ (.A(\i_ca.ca_wr_douta[6] ),
    .B(_1092_),
    .X(_1114_));
 sky130_fd_sc_hd__a221o_1 _2441_ (.A1(\i_ca.hs_write_dbus_wr_data_const[6] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[6] ),
    .C1(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(\i_ca.ca_wr_dina[6] ),
    .A1(_1115_),
    .S(_1097_),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _2443_ (.A(_1116_),
    .X(_0440_));
 sky130_fd_sc_hd__and2_1 _2444_ (.A(\i_ca.ca_wr_douta[7] ),
    .B(_1092_),
    .X(_1117_));
 sky130_fd_sc_hd__a221o_1 _2445_ (.A1(\i_ca.hs_write_dbus_wr_data_const[7] ),
    .A2(_1088_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[7] ),
    .C1(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__mux2_1 _2446_ (.A0(\i_ca.ca_wr_dina[7] ),
    .A1(_1118_),
    .S(_1097_),
    .X(_1119_));
 sky130_fd_sc_hd__clkbuf_1 _2447_ (.A(_1119_),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _2448_ (.A(\i_ca.ca_wr_douta[8] ),
    .B(_1092_),
    .X(_1120_));
 sky130_fd_sc_hd__a221o_1 _2449_ (.A1(\i_ca.hs_write_dbus_wr_data_const[8] ),
    .A2(_1087_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[8] ),
    .C1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(\i_ca.ca_wr_dina[8] ),
    .A1(_1121_),
    .S(_1097_),
    .X(_1122_));
 sky130_fd_sc_hd__clkbuf_1 _2451_ (.A(_1122_),
    .X(_0442_));
 sky130_fd_sc_hd__buf_4 _2452_ (.A(_1087_),
    .X(_1123_));
 sky130_fd_sc_hd__buf_4 _2453_ (.A(_1089_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_4 _2454_ (.A(_1091_),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _2455_ (.A1(\i_ca.ca_insert_time[9] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[9] ),
    .X(_1126_));
 sky130_fd_sc_hd__a21o_1 _2456_ (.A1(\i_ca.hs_write_dbus_wr_data_const[9] ),
    .A2(_1123_),
    .B1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(\i_ca.ca_wr_dina[9] ),
    .A1(_1127_),
    .S(_1097_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_1 _2458_ (.A(_1128_),
    .X(_0443_));
 sky130_fd_sc_hd__a22o_1 _2459_ (.A1(\i_ca.ca_insert_time[10] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[10] ),
    .X(_1129_));
 sky130_fd_sc_hd__a21o_1 _2460_ (.A1(\i_ca.hs_write_dbus_wr_data_const[10] ),
    .A2(_1123_),
    .B1(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__buf_4 _2461_ (.A(_1096_),
    .X(_1131_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(\i_ca.ca_wr_dina[10] ),
    .A1(_1130_),
    .S(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _2463_ (.A(_1132_),
    .X(_0444_));
 sky130_fd_sc_hd__a22o_1 _2464_ (.A1(\i_ca.ca_insert_time[11] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[11] ),
    .X(_1133_));
 sky130_fd_sc_hd__a21o_1 _2465_ (.A1(\i_ca.hs_write_dbus_wr_data_const[11] ),
    .A2(_1123_),
    .B1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(\i_ca.ca_wr_dina[11] ),
    .A1(_1134_),
    .S(_1131_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _2467_ (.A(_1135_),
    .X(_0445_));
 sky130_fd_sc_hd__a22o_1 _2468_ (.A1(\i_ca.ca_insert_time[12] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[12] ),
    .X(_1136_));
 sky130_fd_sc_hd__a21o_1 _2469_ (.A1(\i_ca.hs_write_dbus_wr_data_const[12] ),
    .A2(_1123_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _2470_ (.A0(\i_ca.ca_wr_dina[12] ),
    .A1(_1137_),
    .S(_1131_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_1 _2471_ (.A(_1138_),
    .X(_0446_));
 sky130_fd_sc_hd__and2_1 _2472_ (.A(\i_ca.ca_wr_douta[13] ),
    .B(_1091_),
    .X(_1139_));
 sky130_fd_sc_hd__a221o_2 _2473_ (.A1(\i_ca.hs_write_dbus_wr_data_const[13] ),
    .A2(_1087_),
    .B1(_1090_),
    .B2(\i_ca.ca_insert_time[13] ),
    .C1(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(\i_ca.ca_wr_dina[13] ),
    .A1(_1140_),
    .S(_1131_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2475_ (.A(_1141_),
    .X(_0447_));
 sky130_fd_sc_hd__and2_1 _2476_ (.A(\i_ca.ca_wr_douta[14] ),
    .B(_1091_),
    .X(_1142_));
 sky130_fd_sc_hd__a221o_1 _2477_ (.A1(\i_ca.hs_write_dbus_wr_data_const[14] ),
    .A2(_1087_),
    .B1(_1124_),
    .B2(\i_ca.ca_insert_time[14] ),
    .C1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(\i_ca.ca_wr_dina[14] ),
    .A1(_1143_),
    .S(_1131_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2479_ (.A(_1144_),
    .X(_0448_));
 sky130_fd_sc_hd__a22o_1 _2480_ (.A1(\i_ca.ca_insert_time[15] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[15] ),
    .X(_1145_));
 sky130_fd_sc_hd__a21o_1 _2481_ (.A1(\i_ca.hs_write_dbus_wr_data_const[15] ),
    .A2(_1123_),
    .B1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(\i_ca.ca_wr_dina[15] ),
    .A1(_1146_),
    .S(_1131_),
    .X(_1147_));
 sky130_fd_sc_hd__clkbuf_1 _2483_ (.A(_1147_),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _2484_ (.A1(\i_ca.ca_insert_time[16] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[16] ),
    .X(_1148_));
 sky130_fd_sc_hd__a21o_1 _2485_ (.A1(\i_ca.hs_write_dbus_wr_data_const[16] ),
    .A2(_1123_),
    .B1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _2486_ (.A0(\i_ca.ca_wr_dina[16] ),
    .A1(_1149_),
    .S(_1131_),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2487_ (.A(_1150_),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _2488_ (.A1(\i_ca.ca_insert_time[17] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[17] ),
    .X(_1151_));
 sky130_fd_sc_hd__a21o_1 _2489_ (.A1(\i_ca.hs_write_dbus_wr_data_const[17] ),
    .A2(_1123_),
    .B1(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(\i_ca.ca_wr_dina[17] ),
    .A1(_1152_),
    .S(_1131_),
    .X(_1153_));
 sky130_fd_sc_hd__clkbuf_1 _2491_ (.A(_1153_),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _2492_ (.A1(\i_ca.ca_insert_time[18] ),
    .A2(_1124_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[18] ),
    .X(_1154_));
 sky130_fd_sc_hd__a21o_1 _2493_ (.A1(\i_ca.hs_write_dbus_wr_data_const[18] ),
    .A2(_1123_),
    .B1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(\i_ca.ca_wr_dina[18] ),
    .A1(_1155_),
    .S(_1131_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2495_ (.A(_1156_),
    .X(_0452_));
 sky130_fd_sc_hd__and2_1 _2496_ (.A(\i_ca.ca_wr_douta[19] ),
    .B(_1091_),
    .X(_1157_));
 sky130_fd_sc_hd__a221o_2 _2497_ (.A1(\i_ca.hs_write_dbus_wr_data_const[19] ),
    .A2(_1087_),
    .B1(_1124_),
    .B2(\i_ca.ca_insert_time[19] ),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(\i_ca.ca_wr_dina[19] ),
    .A1(_1158_),
    .S(_1131_),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _2499_ (.A(_1159_),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _2500_ (.A1(\i_ca.ca_insert_time[20] ),
    .A2(_1089_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[20] ),
    .X(_1160_));
 sky130_fd_sc_hd__a21o_1 _2501_ (.A1(\i_ca.hs_write_dbus_wr_data_const[20] ),
    .A2(_1123_),
    .B1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(\i_ca.ca_wr_dina[20] ),
    .A1(_1161_),
    .S(_1096_),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _2503_ (.A(_1162_),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _2504_ (.A1(\i_ca.ca_insert_time[21] ),
    .A2(_1089_),
    .B1(_1125_),
    .B2(\i_ca.ca_wr_douta[21] ),
    .X(_1163_));
 sky130_fd_sc_hd__a21o_1 _2505_ (.A1(\i_ca.hs_write_dbus_wr_data_const[21] ),
    .A2(_1088_),
    .B1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(\i_ca.ca_wr_dina[21] ),
    .A1(_1164_),
    .S(_1096_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_1165_),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _2508_ (.A1(\i_ca.ca_insert_time[22] ),
    .A2(_1089_),
    .B1(_1092_),
    .B2(\i_ca.ca_wr_douta[22] ),
    .X(_1166_));
 sky130_fd_sc_hd__a21o_1 _2509_ (.A1(\i_ca.hs_write_dbus_wr_data_const[22] ),
    .A2(_1088_),
    .B1(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(\i_ca.ca_wr_dina[22] ),
    .A1(_1167_),
    .S(_1096_),
    .X(_1168_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_1168_),
    .X(_0456_));
 sky130_fd_sc_hd__a211o_1 _2512_ (.A1(\i_ca.ca_wr_douta[32] ),
    .A2(_0790_),
    .B1(\i_ca.ca_wr_fsm_state[15] ),
    .C1(_1034_),
    .X(_1169_));
 sky130_fd_sc_hd__a21o_1 _2513_ (.A1(\i_ca.ca_wr_sync_update ),
    .A2(_0788_),
    .B1(_0705_),
    .X(_1170_));
 sky130_fd_sc_hd__and3_1 _2514_ (.A(_0858_),
    .B(_1095_),
    .C(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(\i_ca.ca_wr_dina[32] ),
    .A1(_1169_),
    .S(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _2516_ (.A(_1172_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(net34),
    .A1(\i_ca.hs_write_tid_wr0_const[0] ),
    .S(_0846_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2518_ (.A(_1173_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(net35),
    .A1(\i_ca.hs_write_tid_wr0_const[1] ),
    .S(_0846_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2520_ (.A(_1174_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(net36),
    .A1(\i_ca.hs_write_tid_wr0_const[2] ),
    .S(_0846_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _2522_ (.A(_1175_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(net2),
    .A1(\i_ca.hs_write_dbus_wr_data_const[0] ),
    .S(_0846_),
    .X(_1176_));
 sky130_fd_sc_hd__clkbuf_1 _2524_ (.A(_1176_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(net13),
    .A1(\i_ca.hs_write_dbus_wr_data_const[1] ),
    .S(_0846_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(_1177_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(net24),
    .A1(\i_ca.hs_write_dbus_wr_data_const[2] ),
    .S(_0846_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(_1178_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(net27),
    .A1(\i_ca.hs_write_dbus_wr_data_const[3] ),
    .S(_0846_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2530_ (.A(_1179_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(net28),
    .A1(\i_ca.hs_write_dbus_wr_data_const[4] ),
    .S(_0846_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(_1180_),
    .X(_0465_));
 sky130_fd_sc_hd__buf_4 _2533_ (.A(_0845_),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(net29),
    .A1(\i_ca.hs_write_dbus_wr_data_const[5] ),
    .S(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__clkbuf_1 _2535_ (.A(_1182_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(net30),
    .A1(\i_ca.hs_write_dbus_wr_data_const[6] ),
    .S(_1181_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _2537_ (.A(_1183_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(net31),
    .A1(\i_ca.hs_write_dbus_wr_data_const[7] ),
    .S(_1181_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2539_ (.A(_1184_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(net32),
    .A1(\i_ca.hs_write_dbus_wr_data_const[8] ),
    .S(_1181_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2541_ (.A(_1185_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(net33),
    .A1(\i_ca.hs_write_dbus_wr_data_const[9] ),
    .S(_1181_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _2543_ (.A(_1186_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(net3),
    .A1(\i_ca.hs_write_dbus_wr_data_const[10] ),
    .S(_1181_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _2545_ (.A(_1187_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(net4),
    .A1(\i_ca.hs_write_dbus_wr_data_const[11] ),
    .S(_1181_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_1188_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(net5),
    .A1(\i_ca.hs_write_dbus_wr_data_const[12] ),
    .S(_1181_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_1189_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(net6),
    .A1(\i_ca.hs_write_dbus_wr_data_const[13] ),
    .S(_1181_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2551_ (.A(_1190_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(net7),
    .A1(\i_ca.hs_write_dbus_wr_data_const[14] ),
    .S(_1181_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2553_ (.A(_1191_),
    .X(_0475_));
 sky130_fd_sc_hd__buf_4 _2554_ (.A(_0845_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(net8),
    .A1(\i_ca.hs_write_dbus_wr_data_const[15] ),
    .S(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_1193_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(net9),
    .A1(\i_ca.hs_write_dbus_wr_data_const[16] ),
    .S(_1192_),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_1194_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(net10),
    .A1(\i_ca.hs_write_dbus_wr_data_const[17] ),
    .S(_1192_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2560_ (.A(_1195_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(net11),
    .A1(\i_ca.hs_write_dbus_wr_data_const[18] ),
    .S(_1192_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_1196_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _2563_ (.A0(net12),
    .A1(\i_ca.hs_write_dbus_wr_data_const[19] ),
    .S(_1192_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_1197_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(net14),
    .A1(\i_ca.hs_write_dbus_wr_data_const[20] ),
    .S(_1192_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(_1198_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(net15),
    .A1(\i_ca.hs_write_dbus_wr_data_const[21] ),
    .S(_1192_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(_1199_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(net16),
    .A1(\i_ca.hs_write_dbus_wr_data_const[22] ),
    .S(_1192_),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_1 _2570_ (.A(_1200_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net17),
    .A1(\i_ca.hs_write_dbus_wr_data_const[23] ),
    .S(_1192_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2572_ (.A(_1201_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net18),
    .A1(\i_ca.hs_write_dbus_wr_data_const[24] ),
    .S(_1192_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2574_ (.A(_1202_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(net19),
    .A1(\i_ca.hs_write_dbus_wr_data_const[25] ),
    .S(_0845_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2576_ (.A(_1203_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _2577_ (.A0(net20),
    .A1(\i_ca.hs_write_dbus_wr_data_const[26] ),
    .S(_0845_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2578_ (.A(_1204_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net21),
    .A1(\i_ca.hs_write_dbus_wr_data_const[27] ),
    .S(_0845_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2580_ (.A(_1205_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(net22),
    .A1(\i_ca.hs_write_dbus_wr_data_const[28] ),
    .S(_0845_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2582_ (.A(_1206_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(net23),
    .A1(\i_ca.hs_write_dbus_wr_data_const[29] ),
    .S(_0845_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2584_ (.A(_1207_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(net25),
    .A1(\i_ca.hs_write_dbus_wr_data_const[30] ),
    .S(_0845_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2586_ (.A(_1208_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(net26),
    .A1(\i_ca.hs_write_dbus_wr_data_const[31] ),
    .S(_0845_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2588_ (.A(_1209_),
    .X(_0492_));
 sky130_fd_sc_hd__inv_2 _2589_ (.A(\i_ca.hs_state_write_const[3] ),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _2590_ (.A(\i_ca.hs_state_write_const[3] ),
    .B(_0846_),
    .Y(_1211_));
 sky130_fd_sc_hd__o32a_1 _2591_ (.A1(_1210_),
    .A2(\i_ca.ca_dbus_valid_meta ),
    .A3(_0766_),
    .B1(_1211_),
    .B2(net306),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(\i_ca.ca_wr_sync_update_done ),
    .A1(\i_ca.ca_wr_sync_update ),
    .S(\i_ca.ca_wr_fsm_state[14] ),
    .X(_1212_));
 sky130_fd_sc_hd__clkbuf_1 _2593_ (.A(_1212_),
    .X(_0494_));
 sky130_fd_sc_hd__and3_1 _2594_ (.A(_0708_),
    .B(_1031_),
    .C(_1033_),
    .X(_1213_));
 sky130_fd_sc_hd__o2bb2a_1 _2595_ (.A1_N(\i_ca.ca_wr_fsm_state[12] ),
    .A2_N(_1031_),
    .B1(_1213_),
    .B2(\i_ca.ca_update_rd_add ),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(\i_ca.ca_insert_time[0] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[0] ),
    .S(_0012_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _2597_ (.A(_1214_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(\i_ca.ca_insert_time[1] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[1] ),
    .S(_0012_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2599_ (.A(_1215_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(\i_ca.ca_insert_time[2] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[2] ),
    .S(_0012_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _2601_ (.A(_1216_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(\i_ca.ca_insert_time[3] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[3] ),
    .S(_0012_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _2603_ (.A(_1217_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(\i_ca.ca_insert_time[4] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[4] ),
    .S(_0012_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _2605_ (.A(_1218_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(\i_ca.ca_insert_time[5] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[5] ),
    .S(_0012_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _2607_ (.A(_1219_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(\i_ca.ca_insert_time[6] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[6] ),
    .S(_0012_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _2609_ (.A(_1220_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(\i_ca.ca_insert_time[7] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[7] ),
    .S(_0012_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2611_ (.A(_1221_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(\i_ca.ca_insert_time[8] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[8] ),
    .S(_0012_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2613_ (.A(_1222_),
    .X(_0504_));
 sky130_fd_sc_hd__buf_6 _2614_ (.A(_0857_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\i_ca.ca_insert_time[9] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[9] ),
    .S(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(_1224_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(\i_ca.ca_insert_time[10] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[10] ),
    .S(_1223_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _2618_ (.A(_1225_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(\i_ca.ca_insert_time[11] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[11] ),
    .S(_1223_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(_1226_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(\i_ca.ca_insert_time[12] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[12] ),
    .S(_1223_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2622_ (.A(_1227_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(\i_ca.ca_insert_time[13] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[13] ),
    .S(_1223_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(_1228_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(\i_ca.ca_insert_time[14] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[14] ),
    .S(_1223_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_1229_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(\i_ca.ca_insert_time[15] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[15] ),
    .S(_1223_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_1230_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(\i_ca.ca_insert_time[16] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[16] ),
    .S(_1223_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2630_ (.A(_1231_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\i_ca.ca_insert_time[17] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[17] ),
    .S(_1223_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2632_ (.A(_1232_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _2633_ (.A0(\i_ca.ca_insert_time[18] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[18] ),
    .S(_1223_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2634_ (.A(_1233_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _2635_ (.A0(\i_ca.ca_insert_time[19] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[19] ),
    .S(_0857_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2636_ (.A(_1234_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(\i_ca.ca_insert_time[20] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[20] ),
    .S(_0857_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _2638_ (.A(_1235_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\i_ca.ca_insert_time[21] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[21] ),
    .S(_0857_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _2640_ (.A(_1236_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(\i_ca.ca_insert_time[22] ),
    .A1(\i_ca.hs_write_dbus_wr_data_const[22] ),
    .S(_0857_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2642_ (.A(_1237_),
    .X(_0518_));
 sky130_fd_sc_hd__a21o_1 _2643_ (.A1(_0718_),
    .A2(_0788_),
    .B1(_0705_),
    .X(_1238_));
 sky130_fd_sc_hd__nor3_1 _2644_ (.A(_0719_),
    .B(\i_ca.ca_wr_fsm_state[1] ),
    .C(\i_ca.ca_wr_fsm_state[0] ),
    .Y(_1239_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_1239_),
    .A1(\i_ca.ca_wr_sync_update ),
    .S(\i_ca.ca_wr_fsm_state[14] ),
    .X(_1240_));
 sky130_fd_sc_hd__a211o_1 _2646_ (.A1(\i_ca.ca_wr_fsm_state[1] ),
    .A2(\i_ca.ca_wr_douta[32] ),
    .B1(_0010_),
    .C1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(_1238_),
    .A1(\i_ca.ca_ready ),
    .S(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1242_),
    .X(_0519_));
 sky130_fd_sc_hd__a21oi_4 _2649_ (.A1(\i_ca.ca_end_of_wr_list ),
    .A2(_0768_),
    .B1(_0841_),
    .Y(_1243_));
 sky130_fd_sc_hd__and2_4 _2650_ (.A(\i_ca.ca_wr_com_const ),
    .B(_1087_),
    .X(_1244_));
 sky130_fd_sc_hd__or2_4 _2651_ (.A(\i_ca.ca_wr_fsm_state[4] ),
    .B(_0001_),
    .X(_1245_));
 sky130_fd_sc_hd__a22o_1 _2652_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[23] ),
    .B1(\i_ca.ca_wr_add_ptr[0] ),
    .B2(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__a221o_1 _2653_ (.A1(\i_ca.ca_wr_add_start[0] ),
    .A2(_1243_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[23] ),
    .C1(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__nand3b_4 _2654_ (.A_N(_0011_),
    .B(_1095_),
    .C(_1170_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(_1247_),
    .A1(\i_ca.ca_wr_dina[23] ),
    .S(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2656_ (.A(_1249_),
    .X(_0520_));
 sky130_fd_sc_hd__clkinv_4 _2657_ (.A(_1248_),
    .Y(_1250_));
 sky130_fd_sc_hd__buf_4 _2658_ (.A(_1243_),
    .X(_1251_));
 sky130_fd_sc_hd__a22o_1 _2659_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[24] ),
    .B1(\i_ca.ca_wr_add_ptr[1] ),
    .B2(_1245_),
    .X(_1252_));
 sky130_fd_sc_hd__a221o_1 _2660_ (.A1(_1070_),
    .A2(_1251_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[24] ),
    .C1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__a211o_1 _2661_ (.A1(\i_ca.ca_wr_add_fill[1] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__o21a_1 _2662_ (.A1(\i_ca.ca_wr_dina[24] ),
    .A2(_1250_),
    .B1(_1254_),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _2663_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[25] ),
    .B1(\i_ca.ca_wr_add_ptr[2] ),
    .B2(_1245_),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _2664_ (.A1(\i_ca.ca_wr_add_start[2] ),
    .A2(_1251_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[25] ),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a211o_1 _2665_ (.A1(\i_ca.ca_wr_add_fill[2] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__o21a_1 _2666_ (.A1(\i_ca.ca_wr_dina[25] ),
    .A2(_1250_),
    .B1(_1257_),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _2667_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[26] ),
    .B1(\i_ca.ca_wr_add_ptr[3] ),
    .B2(_1245_),
    .X(_1258_));
 sky130_fd_sc_hd__a221o_1 _2668_ (.A1(\i_ca.ca_wr_add_start[3] ),
    .A2(_1251_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[26] ),
    .C1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a211o_1 _2669_ (.A1(\i_ca.ca_wr_add_fill[3] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__o21a_1 _2670_ (.A1(\i_ca.ca_wr_dina[26] ),
    .A2(_1250_),
    .B1(_1260_),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _2671_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[27] ),
    .B1(\i_ca.ca_wr_add_ptr[4] ),
    .B2(_1245_),
    .X(_1261_));
 sky130_fd_sc_hd__a221o_1 _2672_ (.A1(\i_ca.ca_wr_add_start[4] ),
    .A2(_1243_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[27] ),
    .C1(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__a211o_1 _2673_ (.A1(\i_ca.ca_wr_add_fill[4] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__o21a_1 _2674_ (.A1(\i_ca.ca_wr_dina[27] ),
    .A2(_1250_),
    .B1(_1263_),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _2675_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[28] ),
    .B1(\i_ca.ca_wr_add_ptr[5] ),
    .B2(_1245_),
    .X(_1264_));
 sky130_fd_sc_hd__a221o_1 _2676_ (.A1(\i_ca.ca_wr_add_start[5] ),
    .A2(_1243_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[28] ),
    .C1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__a211o_1 _2677_ (.A1(\i_ca.ca_wr_add_fill[5] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__o21a_1 _2678_ (.A1(\i_ca.ca_wr_dina[28] ),
    .A2(_1250_),
    .B1(_1266_),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _2679_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[29] ),
    .B1(\i_ca.ca_wr_add_ptr[6] ),
    .B2(_1245_),
    .X(_1267_));
 sky130_fd_sc_hd__a221o_1 _2680_ (.A1(\i_ca.ca_wr_add_start[6] ),
    .A2(_1243_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[29] ),
    .C1(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__a211o_1 _2681_ (.A1(\i_ca.ca_wr_add_fill[6] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__o21a_1 _2682_ (.A1(\i_ca.ca_wr_dina[29] ),
    .A2(_1250_),
    .B1(_1269_),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _2683_ (.A1(_0790_),
    .A2(\i_ca.ca_wr_douta[30] ),
    .B1(\i_ca.ca_wr_add_ptr[7] ),
    .B2(_1245_),
    .X(_1270_));
 sky130_fd_sc_hd__a221o_1 _2684_ (.A1(\i_ca.ca_wr_add_start[7] ),
    .A2(_1243_),
    .B1(_1244_),
    .B2(\i_ca.hs_write_dbus_wr_data_const[30] ),
    .C1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a211o_1 _2685_ (.A1(\i_ca.ca_wr_add_fill[7] ),
    .A2(_0025_),
    .B1(_1248_),
    .C1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__o21a_1 _2686_ (.A1(\i_ca.ca_wr_dina[30] ),
    .A2(_1250_),
    .B1(_1272_),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _2687_ (.A1(\i_ca.ca_wr_add_start[8] ),
    .A2(_1251_),
    .B1(_1245_),
    .B2(\i_ca.ca_wr_add_ptr[8] ),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _2688_ (.A1(\i_ca.ca_wr_add_fill[8] ),
    .A2(_0025_),
    .B1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a31o_1 _2689_ (.A1(\i_ca.ca_wr_com_const ),
    .A2(\i_ca.hs_write_dbus_wr_data_const[31] ),
    .A3(_1123_),
    .B1(_1248_),
    .X(_1275_));
 sky130_fd_sc_hd__o22a_1 _2690_ (.A1(\i_ca.ca_wr_dina[31] ),
    .A2(_1250_),
    .B1(_1274_),
    .B2(_1275_),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _2691_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[0] ),
    .B1(\i_ca.ca_wr_add_start[0] ),
    .B2(_1085_),
    .X(_1276_));
 sky130_fd_sc_hd__o21ai_1 _2692_ (.A1(\i_ca.ca_wr_com_const ),
    .A2(_0788_),
    .B1(_0719_),
    .Y(_1277_));
 sky130_fd_sc_hd__and4bb_1 _2693_ (.A_N(_0711_),
    .B_N(_1243_),
    .C(_1277_),
    .D(_1059_),
    .X(_1278_));
 sky130_fd_sc_hd__buf_6 _2694_ (.A(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(\i_ca.ca_wr_add_ptr[0] ),
    .A1(_1276_),
    .S(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2696_ (.A(_1280_),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_1 _2697_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[1] ),
    .B1(_1070_),
    .B2(_1085_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(\i_ca.ca_wr_add_ptr[1] ),
    .A1(_1281_),
    .S(_1279_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2699_ (.A(_1282_),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _2700_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[2] ),
    .B1(\i_ca.ca_wr_add_start[2] ),
    .B2(_1085_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(\i_ca.ca_wr_add_ptr[2] ),
    .A1(_1283_),
    .S(_1279_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2702_ (.A(_1284_),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _2703_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[3] ),
    .B1(\i_ca.ca_wr_add_start[3] ),
    .B2(_1085_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(\i_ca.ca_wr_add_ptr[3] ),
    .A1(_1285_),
    .S(_1279_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2705_ (.A(_1286_),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _2706_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[4] ),
    .B1(\i_ca.ca_wr_add_start[4] ),
    .B2(_1085_),
    .X(_1287_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(\i_ca.ca_wr_add_ptr[4] ),
    .A1(_1287_),
    .S(_1279_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2708_ (.A(_1288_),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_1 _2709_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[5] ),
    .B1(\i_ca.ca_wr_add_start[5] ),
    .B2(_1085_),
    .X(_1289_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\i_ca.ca_wr_add_ptr[5] ),
    .A1(_1289_),
    .S(_1279_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2711_ (.A(_1290_),
    .X(_0534_));
 sky130_fd_sc_hd__a22o_1 _2712_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[6] ),
    .B1(\i_ca.ca_wr_add_start[6] ),
    .B2(_1085_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(\i_ca.ca_wr_add_ptr[6] ),
    .A1(_1291_),
    .S(_1279_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1292_),
    .X(_0535_));
 sky130_fd_sc_hd__a22o_1 _2715_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[7] ),
    .B1(\i_ca.ca_wr_add_start[7] ),
    .B2(_1085_),
    .X(_1293_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\i_ca.ca_wr_add_ptr[7] ),
    .A1(_1293_),
    .S(_1279_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2717_ (.A(_1294_),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _2718_ (.A1(_1060_),
    .A2(\i_ca.ca_wr_add[8] ),
    .B1(\i_ca.ca_wr_add_start[8] ),
    .B2(_1085_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(\i_ca.ca_wr_add_ptr[8] ),
    .A1(_1295_),
    .S(_1279_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2720_ (.A(_1296_),
    .X(_0537_));
 sky130_fd_sc_hd__o211a_1 _2721_ (.A1(_0720_),
    .A2(_0708_),
    .B1(_0841_),
    .C1(_1277_),
    .X(_0538_));
 sky130_fd_sc_hd__or3_2 _2722_ (.A(\i_ca.ca_wr_fsm_state[4] ),
    .B(\i_ca.ca_wr_fsm_state[3] ),
    .C(\i_ca.ca_wr_fsm_state[12] ),
    .X(_1297_));
 sky130_fd_sc_hd__or3_4 _2723_ (.A(\i_ca.ca_wr_fsm_state[14] ),
    .B(\i_ca.ca_wr_fsm_state[13] ),
    .C(\i_ca.ca_wr_fsm_state[11] ),
    .X(_1298_));
 sky130_fd_sc_hd__nor3_4 _2724_ (.A(_1059_),
    .B(_1297_),
    .C(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__a211o_4 _2725_ (.A1(_0764_),
    .A2(_1299_),
    .B1(_0011_),
    .C1(_0717_),
    .X(_1300_));
 sky130_fd_sc_hd__or2_4 _2726_ (.A(_0707_),
    .B(_1298_),
    .X(_1301_));
 sky130_fd_sc_hd__a31o_1 _2727_ (.A1(\i_ca.ca_wr_fsm_state[7] ),
    .A2(\i_ca.ca_wr_douta[32] ),
    .A3(\i_ca.ca_wr_douta[23] ),
    .B1(\i_ca.ca_wr_fsm_state[3] ),
    .X(_1302_));
 sky130_fd_sc_hd__a311o_1 _2728_ (.A1(_0719_),
    .A2(\i_ca.hs_write_tid_wr0_const[0] ),
    .A3(_1062_),
    .B1(_1299_),
    .C1(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__a221o_1 _2729_ (.A1(\i_ca.ca_wr_add_ptr[0] ),
    .A2(_0787_),
    .B1(_1301_),
    .B2(\i_ca.ca_wr_add_start[0] ),
    .C1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__a31o_1 _2730_ (.A1(_0774_),
    .A2(\i_ca.ca_wr_dina[23] ),
    .A3(_1251_),
    .B1(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__a21oi_1 _2731_ (.A1(\i_ca.ca_wr_add[0] ),
    .A2(_1299_),
    .B1(_1300_),
    .Y(_1306_));
 sky130_fd_sc_hd__a22o_1 _2732_ (.A1(\i_ca.ca_wr_add[0] ),
    .A2(_1300_),
    .B1(_1305_),
    .B2(_1306_),
    .X(_0539_));
 sky130_fd_sc_hd__a22o_1 _2733_ (.A1(\i_ca.ca_wr_douta[24] ),
    .A2(_0001_),
    .B1(_1298_),
    .B2(_1070_),
    .X(_1307_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_1070_),
    .A1(\i_ca.hs_write_tid_wr0_const[1] ),
    .S(_1062_),
    .X(_1308_));
 sky130_fd_sc_hd__or2_4 _2735_ (.A(_0711_),
    .B(_1297_),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(\i_ca.ca_wr_dina[24] ),
    .A1(\i_ca.ca_wr_add_fill[1] ),
    .S(_0708_),
    .X(_1310_));
 sky130_fd_sc_hd__a22o_1 _2737_ (.A1(\i_ca.ca_wr_add_ptr[1] ),
    .A2(_0787_),
    .B1(_1243_),
    .B2(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__a221o_1 _2738_ (.A1(_0720_),
    .A2(_1308_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[1] ),
    .C1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__nand2_1 _2739_ (.A(\i_ca.ca_wr_add[0] ),
    .B(\i_ca.ca_wr_add[1] ),
    .Y(_1313_));
 sky130_fd_sc_hd__or2_1 _2740_ (.A(\i_ca.ca_wr_add[0] ),
    .B(\i_ca.ca_wr_add[1] ),
    .X(_1314_));
 sky130_fd_sc_hd__a31o_1 _2741_ (.A1(_1313_),
    .A2(_1299_),
    .A3(_1314_),
    .B1(_1300_),
    .X(_1315_));
 sky130_fd_sc_hd__or3_4 _2742_ (.A(_1059_),
    .B(_1297_),
    .C(_1298_),
    .X(_1316_));
 sky130_fd_sc_hd__o221a_4 _2743_ (.A1(\i_ca.ca_end_of_wr_list ),
    .A2(_0858_),
    .B1(_1316_),
    .B2(\i_ca.ca_wr_fsm_state[0] ),
    .C1(_1065_),
    .X(_1317_));
 sky130_fd_sc_hd__o32a_1 _2744_ (.A1(_1307_),
    .A2(_1312_),
    .A3(_1315_),
    .B1(_1317_),
    .B2(\i_ca.ca_wr_add[1] ),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _2745_ (.A(_0712_),
    .Y(_1318_));
 sky130_fd_sc_hd__a21o_1 _2746_ (.A1(\i_ca.ca_wr_add[0] ),
    .A2(\i_ca.ca_wr_add[1] ),
    .B1(\i_ca.ca_wr_add[2] ),
    .X(_1319_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(\i_ca.ca_wr_add_start[2] ),
    .A1(\i_ca.hs_write_tid_wr0_const[2] ),
    .S(_1062_),
    .X(_1320_));
 sky130_fd_sc_hd__a22o_1 _2748_ (.A1(\i_ca.ca_wr_add_fill[2] ),
    .A2(_1309_),
    .B1(_1320_),
    .B2(_0719_),
    .X(_1321_));
 sky130_fd_sc_hd__a221o_1 _2749_ (.A1(\i_ca.ca_wr_douta[25] ),
    .A2(_0001_),
    .B1(_1298_),
    .B2(\i_ca.ca_wr_add_start[2] ),
    .C1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a31o_1 _2750_ (.A1(_1318_),
    .A2(_1299_),
    .A3(_1319_),
    .B1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(\i_ca.ca_wr_dina[25] ),
    .A1(\i_ca.ca_wr_add_fill[2] ),
    .S(_0708_),
    .X(_1324_));
 sky130_fd_sc_hd__a221o_1 _2752_ (.A1(\i_ca.ca_wr_add_ptr[2] ),
    .A2(_0787_),
    .B1(_1251_),
    .B2(_1324_),
    .C1(_1300_),
    .X(_1325_));
 sky130_fd_sc_hd__o22a_1 _2753_ (.A1(\i_ca.ca_wr_add[2] ),
    .A2(_1317_),
    .B1(_1323_),
    .B2(_1325_),
    .X(_0541_));
 sky130_fd_sc_hd__xor2_1 _2754_ (.A(\i_ca.ca_wr_add[3] ),
    .B(_0712_),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(\i_ca.ca_wr_dina[26] ),
    .A1(\i_ca.ca_wr_add_fill[3] ),
    .S(\i_ca.ca_wr_add_start_marker ),
    .X(_1327_));
 sky130_fd_sc_hd__a22o_1 _2756_ (.A1(\i_ca.ca_wr_add_ptr[3] ),
    .A2(_0787_),
    .B1(_1243_),
    .B2(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a221o_1 _2757_ (.A1(\i_ca.ca_wr_douta[26] ),
    .A2(_0001_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[3] ),
    .C1(_1299_),
    .X(_1329_));
 sky130_fd_sc_hd__a211o_1 _2758_ (.A1(\i_ca.ca_wr_add_start[3] ),
    .A2(_1301_),
    .B1(_1328_),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__o211a_1 _2759_ (.A1(_1316_),
    .A2(_1326_),
    .B1(_1330_),
    .C1(_1317_),
    .X(_1331_));
 sky130_fd_sc_hd__a21o_1 _2760_ (.A1(\i_ca.ca_wr_add[3] ),
    .A2(_1300_),
    .B1(_1331_),
    .X(_0542_));
 sky130_fd_sc_hd__a221o_1 _2761_ (.A1(\i_ca.ca_wr_douta[27] ),
    .A2(_0001_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[4] ),
    .C1(_1299_),
    .X(_1332_));
 sky130_fd_sc_hd__mux2_1 _2762_ (.A0(\i_ca.ca_wr_dina[27] ),
    .A1(\i_ca.ca_wr_add_fill[4] ),
    .S(_0708_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_1 _2763_ (.A1(\i_ca.ca_wr_add_ptr[4] ),
    .A2(_0787_),
    .B1(_1251_),
    .B2(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__a211o_1 _2764_ (.A1(\i_ca.ca_wr_add_start[4] ),
    .A2(_1301_),
    .B1(_1332_),
    .C1(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__a21oi_1 _2765_ (.A1(\i_ca.ca_wr_add[3] ),
    .A2(_0712_),
    .B1(\i_ca.ca_wr_add[4] ),
    .Y(_1336_));
 sky130_fd_sc_hd__o211a_1 _2766_ (.A1(_0713_),
    .A2(_1336_),
    .B1(_1299_),
    .C1(_0715_),
    .X(_1337_));
 sky130_fd_sc_hd__nor2_1 _2767_ (.A(_1300_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__a22o_1 _2768_ (.A1(\i_ca.ca_wr_add[4] ),
    .A2(_1300_),
    .B1(_1335_),
    .B2(_1338_),
    .X(_0543_));
 sky130_fd_sc_hd__nor2_1 _2769_ (.A(\i_ca.ca_wr_add[5] ),
    .B(_0713_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21a_1 _2770_ (.A1(_0714_),
    .A2(_1316_),
    .B1(_1317_),
    .X(_1340_));
 sky130_fd_sc_hd__a21oi_1 _2771_ (.A1(_1317_),
    .A2(_1339_),
    .B1(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__a22o_1 _2772_ (.A1(\i_ca.ca_wr_douta[28] ),
    .A2(_0001_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[5] ),
    .X(_1342_));
 sky130_fd_sc_hd__a21o_1 _2773_ (.A1(\i_ca.ca_wr_add_start[5] ),
    .A2(_1301_),
    .B1(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(\i_ca.ca_wr_dina[28] ),
    .A1(\i_ca.ca_wr_add_fill[5] ),
    .S(_0708_),
    .X(_1344_));
 sky130_fd_sc_hd__a22o_1 _2775_ (.A1(\i_ca.ca_wr_add_ptr[5] ),
    .A2(_0787_),
    .B1(_1251_),
    .B2(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__o32a_1 _2776_ (.A1(_1341_),
    .A2(_1343_),
    .A3(_1345_),
    .B1(_1317_),
    .B2(\i_ca.ca_wr_add[5] ),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\i_ca.ca_wr_dina[29] ),
    .A1(\i_ca.ca_wr_add_fill[6] ),
    .S(_0708_),
    .X(_1346_));
 sky130_fd_sc_hd__a22o_1 _2778_ (.A1(\i_ca.ca_wr_douta[29] ),
    .A2(_0001_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[6] ),
    .X(_1347_));
 sky130_fd_sc_hd__a221o_1 _2779_ (.A1(\i_ca.ca_wr_add_start[6] ),
    .A2(_1301_),
    .B1(_1346_),
    .B2(_1251_),
    .C1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a21oi_1 _2780_ (.A1(\i_ca.ca_wr_add_ptr[6] ),
    .A2(_0787_),
    .B1(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__and3_1 _2781_ (.A(\i_ca.ca_wr_add[5] ),
    .B(\i_ca.ca_wr_add[6] ),
    .C(_0713_),
    .X(_1350_));
 sky130_fd_sc_hd__o31a_1 _2782_ (.A1(_0716_),
    .A2(_1316_),
    .A3(_1350_),
    .B1(_1317_),
    .X(_1351_));
 sky130_fd_sc_hd__o2bb2a_1 _2783_ (.A1_N(_1349_),
    .A2_N(_1351_),
    .B1(\i_ca.ca_wr_add[6] ),
    .B2(_1340_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(\i_ca.ca_wr_dina[30] ),
    .A1(\i_ca.ca_wr_add_fill[7] ),
    .S(_0708_),
    .X(_1352_));
 sky130_fd_sc_hd__a22o_1 _2785_ (.A1(\i_ca.ca_wr_douta[30] ),
    .A2(_0001_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[7] ),
    .X(_1353_));
 sky130_fd_sc_hd__a21o_1 _2786_ (.A1(\i_ca.ca_wr_add_start[7] ),
    .A2(_1301_),
    .B1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a221o_1 _2787_ (.A1(\i_ca.ca_wr_add_ptr[7] ),
    .A2(_0787_),
    .B1(_1251_),
    .B2(_1352_),
    .C1(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__nand2_1 _2788_ (.A(\i_ca.ca_wr_add[7] ),
    .B(_1350_),
    .Y(_1356_));
 sky130_fd_sc_hd__a21o_1 _2789_ (.A1(_1299_),
    .A2(_1356_),
    .B1(_1300_),
    .X(_1357_));
 sky130_fd_sc_hd__o31a_1 _2790_ (.A1(\i_ca.ca_wr_add[7] ),
    .A2(_1300_),
    .A3(_1350_),
    .B1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__o22a_1 _2791_ (.A1(\i_ca.ca_wr_add[7] ),
    .A2(_1317_),
    .B1(_1355_),
    .B2(_1358_),
    .X(_0546_));
 sky130_fd_sc_hd__nor3_1 _2792_ (.A(\i_ca.ca_wr_add[8] ),
    .B(_1316_),
    .C(_1356_),
    .Y(_1359_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(\i_ca.ca_wr_dina[31] ),
    .A1(\i_ca.ca_wr_add_fill[8] ),
    .S(\i_ca.ca_wr_add_start_marker ),
    .X(_1360_));
 sky130_fd_sc_hd__and2_1 _2794_ (.A(_1243_),
    .B(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__a221o_1 _2795_ (.A1(\i_ca.ca_wr_add_start[8] ),
    .A2(_1301_),
    .B1(_1309_),
    .B2(\i_ca.ca_wr_add_fill[8] ),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__a211o_1 _2796_ (.A1(\i_ca.ca_wr_add_ptr[8] ),
    .A2(_0787_),
    .B1(_1359_),
    .C1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__a22o_1 _2797_ (.A1(\i_ca.ca_wr_add[8] ),
    .A2(_1357_),
    .B1(_1363_),
    .B2(_1317_),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_1 _2798_ (.A(_0723_),
    .B(\i_ca.ca_rd_fsm_state[6] ),
    .Y(_1364_));
 sky130_fd_sc_hd__a22o_1 _2799_ (.A1(\i_ca.ca_wr_sync_update ),
    .A2(_1364_),
    .B1(_0771_),
    .B2(\i_ca.ca_rd_fsm_state[6] ),
    .X(_0548_));
 sky130_fd_sc_hd__or3_1 _2800_ (.A(\i_ca.ca_update_rd_add ),
    .B(\i_ca.ca_rd_fsm_state[6] ),
    .C(\i_ca.ca_rd_fsm_state[3] ),
    .X(_1365_));
 sky130_fd_sc_hd__buf_4 _2801_ (.A(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(_0773_),
    .A1(_1366_),
    .S(\i_ca.ca_wr_add_start[0] ),
    .X(_1367_));
 sky130_fd_sc_hd__o2bb2a_1 _2803_ (.A1_N(_0773_),
    .A2_N(_0780_),
    .B1(\i_ca.ca_wr_sync_update_done ),
    .B2(_1364_),
    .X(_1368_));
 sky130_fd_sc_hd__o31a_4 _2804_ (.A1(\i_ca.ca_rd_fsm_state[5] ),
    .A2(\i_ca.ca_rd_fsm_state[0] ),
    .A3(_1366_),
    .B1(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\i_ca.ca_rd_add[0] ),
    .A1(_1367_),
    .S(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _2806_ (.A(_1370_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _2807_ (.A(\i_ca.ca_wr_add_start[0] ),
    .B(_1070_),
    .Y(_1371_));
 sky130_fd_sc_hd__or2_1 _2808_ (.A(\i_ca.ca_wr_add_start[0] ),
    .B(_1070_),
    .X(_1372_));
 sky130_fd_sc_hd__a32o_1 _2809_ (.A1(_0773_),
    .A2(_1371_),
    .A3(_1372_),
    .B1(_1366_),
    .B2(_1070_),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(\i_ca.ca_rd_add[1] ),
    .A1(_1373_),
    .S(_1369_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _2811_ (.A(_1374_),
    .X(_0550_));
 sky130_fd_sc_hd__nand3_1 _2812_ (.A(\i_ca.ca_wr_add_start[0] ),
    .B(_1070_),
    .C(\i_ca.ca_wr_add_start[2] ),
    .Y(_1375_));
 sky130_fd_sc_hd__a21o_1 _2813_ (.A1(\i_ca.ca_wr_add_start[0] ),
    .A2(_1070_),
    .B1(\i_ca.ca_wr_add_start[2] ),
    .X(_1376_));
 sky130_fd_sc_hd__a32o_1 _2814_ (.A1(_0773_),
    .A2(_1375_),
    .A3(_1376_),
    .B1(_1366_),
    .B2(\i_ca.ca_wr_add_start[2] ),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(\i_ca.ca_rd_add[2] ),
    .A1(_1377_),
    .S(_1369_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _2816_ (.A(_1378_),
    .X(_0551_));
 sky130_fd_sc_hd__o21bai_1 _2817_ (.A1(\i_ca.ca_update_rd_add ),
    .A2(_1375_),
    .B1_N(\i_ca.ca_wr_add_start[3] ),
    .Y(_1379_));
 sky130_fd_sc_hd__and4_2 _2818_ (.A(\i_ca.ca_wr_add_start[0] ),
    .B(\i_ca.ca_wr_add_start[1] ),
    .C(\i_ca.ca_wr_add_start[2] ),
    .D(\i_ca.ca_wr_add_start[3] ),
    .X(_1380_));
 sky130_fd_sc_hd__inv_2 _2819_ (.A(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__a32o_1 _2820_ (.A1(\i_ca.ca_rd_fsm_state[5] ),
    .A2(_1379_),
    .A3(_1381_),
    .B1(\i_ca.ca_wr_add_start[3] ),
    .B2(_1366_),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(\i_ca.ca_rd_add[3] ),
    .A1(_1382_),
    .S(_1369_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _2822_ (.A(_1383_),
    .X(_0552_));
 sky130_fd_sc_hd__inv_2 _2823_ (.A(_1366_),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _2824_ (.A(_1384_),
    .B(_1380_),
    .Y(_1385_));
 sky130_fd_sc_hd__mux2_1 _2825_ (.A0(_1380_),
    .A1(_1385_),
    .S(\i_ca.ca_wr_add_start[4] ),
    .X(_1386_));
 sky130_fd_sc_hd__o32a_1 _2826_ (.A1(\i_ca.ca_wr_add_start[4] ),
    .A2(_0773_),
    .A3(_1384_),
    .B1(_1386_),
    .B2(_0772_),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(\i_ca.ca_rd_add[4] ),
    .A1(_1387_),
    .S(_1369_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _2828_ (.A(_1388_),
    .X(_0553_));
 sky130_fd_sc_hd__a31o_1 _2829_ (.A1(_0723_),
    .A2(\i_ca.ca_wr_add_start[4] ),
    .A3(_1380_),
    .B1(\i_ca.ca_wr_add_start[5] ),
    .X(_1389_));
 sky130_fd_sc_hd__and3_1 _2830_ (.A(\i_ca.ca_wr_add_start[4] ),
    .B(\i_ca.ca_wr_add_start[5] ),
    .C(_1380_),
    .X(_1390_));
 sky130_fd_sc_hd__inv_2 _2831_ (.A(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a32o_1 _2832_ (.A1(\i_ca.ca_rd_fsm_state[5] ),
    .A2(_1389_),
    .A3(_1391_),
    .B1(\i_ca.ca_wr_add_start[5] ),
    .B2(_1366_),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\i_ca.ca_rd_add[5] ),
    .A1(_1392_),
    .S(_1369_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _2834_ (.A(_1393_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _2835_ (.A(\i_ca.ca_wr_add_start[6] ),
    .B(_1390_),
    .X(_1394_));
 sky130_fd_sc_hd__nand2_1 _2836_ (.A(\i_ca.ca_wr_add_start[6] ),
    .B(_1390_),
    .Y(_1395_));
 sky130_fd_sc_hd__a32o_1 _2837_ (.A1(_0773_),
    .A2(_1394_),
    .A3(_1395_),
    .B1(_1366_),
    .B2(\i_ca.ca_wr_add_start[6] ),
    .X(_1396_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(\i_ca.ca_rd_add[6] ),
    .A1(_1396_),
    .S(_1369_),
    .X(_1397_));
 sky130_fd_sc_hd__clkbuf_1 _2839_ (.A(_1397_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _2840_ (.A(\i_ca.ca_update_rd_add ),
    .B(\i_ca.ca_wr_add_start[7] ),
    .Y(_1398_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(_1398_),
    .A1(\i_ca.ca_wr_add_start[7] ),
    .S(_1395_),
    .X(_1399_));
 sky130_fd_sc_hd__a22o_1 _2842_ (.A1(\i_ca.ca_wr_add_start[7] ),
    .A2(_1366_),
    .B1(_1399_),
    .B2(\i_ca.ca_rd_fsm_state[5] ),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(\i_ca.ca_rd_add[7] ),
    .A1(_1400_),
    .S(_1369_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _2844_ (.A(_1401_),
    .X(_0556_));
 sky130_fd_sc_hd__o21ai_1 _2845_ (.A1(_0726_),
    .A2(_0728_),
    .B1(net307),
    .Y(_1402_));
 sky130_fd_sc_hd__o2bb2a_1 _2846_ (.A1_N(\i_ca.ca_match_hs_state[2] ),
    .A2_N(_1402_),
    .B1(_0005_),
    .B2(net307),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_2 _2847_ (.A(_0727_),
    .B(_0034_),
    .Y(_1403_));
 sky130_fd_sc_hd__buf_4 _2848_ (.A(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(\i_ca.ca_rd_doutb[0] ),
    .A1(net275),
    .S(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1405_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\i_ca.ca_rd_doutb[1] ),
    .A1(net286),
    .S(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _2852_ (.A(_1406_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\i_ca.ca_rd_doutb[2] ),
    .A1(net297),
    .S(_1404_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1407_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\i_ca.ca_rd_doutb[3] ),
    .A1(net299),
    .S(_1404_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _2856_ (.A(_1408_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\i_ca.ca_rd_doutb[4] ),
    .A1(net300),
    .S(_1404_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _2858_ (.A(_1409_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\i_ca.ca_rd_doutb[5] ),
    .A1(net301),
    .S(_1404_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(_1410_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(\i_ca.ca_rd_doutb[6] ),
    .A1(net302),
    .S(_1404_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _2862_ (.A(_1411_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(\i_ca.ca_rd_doutb[7] ),
    .A1(net303),
    .S(_1404_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _2864_ (.A(_1412_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\i_ca.ca_rd_doutb[8] ),
    .A1(net304),
    .S(_1404_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1413_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(\i_ca.ca_rd_doutb[9] ),
    .A1(net305),
    .S(_1404_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _2868_ (.A(_1414_),
    .X(_0567_));
 sky130_fd_sc_hd__buf_4 _2869_ (.A(_1403_),
    .X(_1415_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\i_ca.ca_rd_doutb[10] ),
    .A1(net276),
    .S(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _2871_ (.A(_1416_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\i_ca.ca_rd_doutb[11] ),
    .A1(net277),
    .S(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _2873_ (.A(_1417_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\i_ca.ca_rd_doutb[12] ),
    .A1(net278),
    .S(_1415_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1418_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\i_ca.ca_rd_doutb[13] ),
    .A1(net279),
    .S(_1415_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1419_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(\i_ca.ca_rd_doutb[14] ),
    .A1(net280),
    .S(_1415_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_1420_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(\i_ca.ca_rd_doutb[15] ),
    .A1(net281),
    .S(_1415_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _2881_ (.A(_1421_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(\i_ca.ca_rd_doutb[16] ),
    .A1(net282),
    .S(_1415_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _2883_ (.A(_1422_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(\i_ca.ca_rd_doutb[17] ),
    .A1(net283),
    .S(_1415_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(_1423_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(\i_ca.ca_rd_doutb[18] ),
    .A1(net284),
    .S(_1415_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _2887_ (.A(_1424_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(\i_ca.ca_rd_doutb[19] ),
    .A1(net285),
    .S(_1415_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _2889_ (.A(_1425_),
    .X(_0577_));
 sky130_fd_sc_hd__buf_4 _2890_ (.A(_1403_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(\i_ca.ca_rd_doutb[20] ),
    .A1(net287),
    .S(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1427_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(\i_ca.ca_rd_doutb[21] ),
    .A1(net288),
    .S(_1426_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _2894_ (.A(_1428_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(\i_ca.ca_rd_doutb[22] ),
    .A1(net289),
    .S(_1426_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _2896_ (.A(_1429_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(\i_ca.ca_rd_doutb[23] ),
    .A1(net290),
    .S(_1426_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_1430_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(\i_ca.ca_rd_doutb[24] ),
    .A1(net291),
    .S(_1426_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _2900_ (.A(_1431_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(\i_ca.ca_rd_doutb[25] ),
    .A1(net292),
    .S(_1426_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _2902_ (.A(_1432_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(\i_ca.ca_rd_doutb[26] ),
    .A1(net293),
    .S(_1426_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _2904_ (.A(_1433_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(\i_ca.ca_rd_doutb[27] ),
    .A1(net294),
    .S(_1426_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _2906_ (.A(_1434_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(\i_ca.ca_rd_doutb[28] ),
    .A1(net295),
    .S(_1426_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _2908_ (.A(_1435_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(\i_ca.ca_rd_doutb[29] ),
    .A1(net296),
    .S(_1426_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1436_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(\i_ca.ca_rd_doutb[30] ),
    .A1(net298),
    .S(_1403_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1437_),
    .X(_0588_));
 sky130_fd_sc_hd__dfrtp_1 _2913_ (.CLK(net754),
    .D(\i_ca.cubev_ca_wea ),
    .RESET_B(_0072_),
    .Q(net382));
 sky130_fd_sc_hd__dfrtp_1 _2914_ (.CLK(net755),
    .D(\i_ca.ca_wr_add[0] ),
    .RESET_B(_0074_),
    .Q(net332));
 sky130_fd_sc_hd__dfrtp_1 _2915_ (.CLK(net756),
    .D(\i_ca.ca_wr_add[1] ),
    .RESET_B(_0076_),
    .Q(net333));
 sky130_fd_sc_hd__dfrtp_1 _2916_ (.CLK(net757),
    .D(\i_ca.ca_wr_add[2] ),
    .RESET_B(_0078_),
    .Q(net334));
 sky130_fd_sc_hd__dfrtp_1 _2917_ (.CLK(net758),
    .D(\i_ca.ca_wr_add[3] ),
    .RESET_B(_0080_),
    .Q(net335));
 sky130_fd_sc_hd__dfrtp_1 _2918_ (.CLK(net759),
    .D(\i_ca.ca_wr_add[4] ),
    .RESET_B(_0082_),
    .Q(net336));
 sky130_fd_sc_hd__dfrtp_1 _2919_ (.CLK(net760),
    .D(\i_ca.ca_wr_add[5] ),
    .RESET_B(_0084_),
    .Q(net337));
 sky130_fd_sc_hd__dfrtp_1 _2920_ (.CLK(net761),
    .D(\i_ca.ca_wr_add[6] ),
    .RESET_B(_0086_),
    .Q(net338));
 sky130_fd_sc_hd__dfrtp_1 _2921_ (.CLK(net762),
    .D(\i_ca.ca_wr_add[7] ),
    .RESET_B(_0088_),
    .Q(net339));
 sky130_fd_sc_hd__dfrtp_1 _2922_ (.CLK(net763),
    .D(\i_ca.ca_wr_dina[0] ),
    .RESET_B(_0090_),
    .Q(net350));
 sky130_fd_sc_hd__dfrtp_1 _2923_ (.CLK(net764),
    .D(\i_ca.ca_wr_dina[1] ),
    .RESET_B(_0092_),
    .Q(net361));
 sky130_fd_sc_hd__dfrtp_1 _2924_ (.CLK(net765),
    .D(\i_ca.ca_wr_dina[2] ),
    .RESET_B(_0094_),
    .Q(net372));
 sky130_fd_sc_hd__dfrtp_1 _2925_ (.CLK(net766),
    .D(\i_ca.ca_wr_dina[3] ),
    .RESET_B(_0096_),
    .Q(net375));
 sky130_fd_sc_hd__dfrtp_1 _2926_ (.CLK(net767),
    .D(\i_ca.ca_wr_dina[4] ),
    .RESET_B(_0098_),
    .Q(net376));
 sky130_fd_sc_hd__dfrtp_1 _2927_ (.CLK(net768),
    .D(\i_ca.ca_wr_dina[5] ),
    .RESET_B(_0100_),
    .Q(net377));
 sky130_fd_sc_hd__dfrtp_1 _2928_ (.CLK(net769),
    .D(\i_ca.ca_wr_dina[6] ),
    .RESET_B(_0102_),
    .Q(net378));
 sky130_fd_sc_hd__dfrtp_1 _2929_ (.CLK(net770),
    .D(\i_ca.ca_wr_dina[7] ),
    .RESET_B(_0104_),
    .Q(net379));
 sky130_fd_sc_hd__dfrtp_1 _2930_ (.CLK(net771),
    .D(\i_ca.ca_wr_dina[8] ),
    .RESET_B(_0106_),
    .Q(net380));
 sky130_fd_sc_hd__dfrtp_1 _2931_ (.CLK(net772),
    .D(\i_ca.ca_wr_dina[9] ),
    .RESET_B(_0108_),
    .Q(net381));
 sky130_fd_sc_hd__dfrtp_1 _2932_ (.CLK(net773),
    .D(\i_ca.ca_wr_dina[10] ),
    .RESET_B(_0110_),
    .Q(net351));
 sky130_fd_sc_hd__dfrtp_1 _2933_ (.CLK(net774),
    .D(\i_ca.ca_wr_dina[11] ),
    .RESET_B(_0112_),
    .Q(net352));
 sky130_fd_sc_hd__dfrtp_1 _2934_ (.CLK(net775),
    .D(\i_ca.ca_wr_dina[12] ),
    .RESET_B(_0114_),
    .Q(net353));
 sky130_fd_sc_hd__dfrtp_1 _2935_ (.CLK(net776),
    .D(\i_ca.ca_wr_dina[13] ),
    .RESET_B(_0116_),
    .Q(net354));
 sky130_fd_sc_hd__dfrtp_1 _2936_ (.CLK(net777),
    .D(\i_ca.ca_wr_dina[14] ),
    .RESET_B(_0118_),
    .Q(net355));
 sky130_fd_sc_hd__dfrtp_1 _2937_ (.CLK(net778),
    .D(\i_ca.ca_wr_dina[15] ),
    .RESET_B(_0120_),
    .Q(net356));
 sky130_fd_sc_hd__dfrtp_1 _2938_ (.CLK(net779),
    .D(\i_ca.ca_wr_dina[16] ),
    .RESET_B(_0122_),
    .Q(net357));
 sky130_fd_sc_hd__dfrtp_1 _2939_ (.CLK(net780),
    .D(\i_ca.ca_wr_dina[17] ),
    .RESET_B(_0124_),
    .Q(net358));
 sky130_fd_sc_hd__dfrtp_1 _2940_ (.CLK(net781),
    .D(\i_ca.ca_wr_dina[18] ),
    .RESET_B(_0126_),
    .Q(net359));
 sky130_fd_sc_hd__dfrtp_1 _2941_ (.CLK(net782),
    .D(\i_ca.ca_wr_dina[19] ),
    .RESET_B(_0128_),
    .Q(net360));
 sky130_fd_sc_hd__dfrtp_1 _2942_ (.CLK(net783),
    .D(\i_ca.ca_wr_dina[20] ),
    .RESET_B(_0130_),
    .Q(net362));
 sky130_fd_sc_hd__dfrtp_1 _2943_ (.CLK(net784),
    .D(\i_ca.ca_wr_dina[21] ),
    .RESET_B(_0132_),
    .Q(net363));
 sky130_fd_sc_hd__dfrtp_1 _2944_ (.CLK(net785),
    .D(\i_ca.ca_wr_dina[22] ),
    .RESET_B(_0134_),
    .Q(net364));
 sky130_fd_sc_hd__dfrtp_1 _2945_ (.CLK(net786),
    .D(\i_ca.ca_wr_dina[23] ),
    .RESET_B(_0136_),
    .Q(net365));
 sky130_fd_sc_hd__dfrtp_1 _2946_ (.CLK(net787),
    .D(\i_ca.ca_wr_dina[24] ),
    .RESET_B(_0138_),
    .Q(net366));
 sky130_fd_sc_hd__dfrtp_1 _2947_ (.CLK(net788),
    .D(\i_ca.ca_wr_dina[25] ),
    .RESET_B(_0140_),
    .Q(net367));
 sky130_fd_sc_hd__dfrtp_1 _2948_ (.CLK(net789),
    .D(\i_ca.ca_wr_dina[26] ),
    .RESET_B(_0142_),
    .Q(net368));
 sky130_fd_sc_hd__dfrtp_1 _2949_ (.CLK(net790),
    .D(\i_ca.ca_wr_dina[27] ),
    .RESET_B(_0144_),
    .Q(net369));
 sky130_fd_sc_hd__dfrtp_1 _2950_ (.CLK(net791),
    .D(\i_ca.ca_wr_dina[28] ),
    .RESET_B(_0146_),
    .Q(net370));
 sky130_fd_sc_hd__dfrtp_1 _2951_ (.CLK(net792),
    .D(\i_ca.ca_wr_dina[29] ),
    .RESET_B(_0148_),
    .Q(net371));
 sky130_fd_sc_hd__dfrtp_1 _2952_ (.CLK(net793),
    .D(\i_ca.ca_wr_dina[30] ),
    .RESET_B(_0150_),
    .Q(net373));
 sky130_fd_sc_hd__dfrtp_1 _2953_ (.CLK(net794),
    .D(\i_ca.ca_wr_dina[32] ),
    .RESET_B(_0152_),
    .Q(net374));
 sky130_fd_sc_hd__dfrtp_1 _2954_ (.CLK(net795),
    .D(\i_ca.ca_rd_add[0] ),
    .RESET_B(_0154_),
    .Q(net340));
 sky130_fd_sc_hd__dfrtp_1 _2955_ (.CLK(net796),
    .D(\i_ca.ca_rd_add[1] ),
    .RESET_B(_0156_),
    .Q(net341));
 sky130_fd_sc_hd__dfrtp_1 _2956_ (.CLK(net797),
    .D(\i_ca.ca_rd_add[2] ),
    .RESET_B(_0158_),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_1 _2957_ (.CLK(net798),
    .D(\i_ca.ca_rd_add[3] ),
    .RESET_B(_0160_),
    .Q(net343));
 sky130_fd_sc_hd__dfrtp_1 _2958_ (.CLK(net799),
    .D(\i_ca.ca_rd_add[4] ),
    .RESET_B(_0162_),
    .Q(net344));
 sky130_fd_sc_hd__dfrtp_1 _2959_ (.CLK(net800),
    .D(\i_ca.ca_rd_add[5] ),
    .RESET_B(_0164_),
    .Q(net345));
 sky130_fd_sc_hd__dfrtp_1 _2960_ (.CLK(net801),
    .D(\i_ca.ca_rd_add[6] ),
    .RESET_B(_0166_),
    .Q(net346));
 sky130_fd_sc_hd__dfrtp_1 _2961_ (.CLK(net802),
    .D(\i_ca.ca_rd_add[7] ),
    .RESET_B(_0168_),
    .Q(net347));
 sky130_fd_sc_hd__dfxtp_2 _2962_ (.CLK(net803),
    .D(net307),
    .Q(net557));
 sky130_fd_sc_hd__dfxtp_1 _2963_ (.CLK(net804),
    .D(net275),
    .Q(net558));
 sky130_fd_sc_hd__dfxtp_1 _2964_ (.CLK(net805),
    .D(net286),
    .Q(net559));
 sky130_fd_sc_hd__dfxtp_1 _2965_ (.CLK(net806),
    .D(net297),
    .Q(net560));
 sky130_fd_sc_hd__dfxtp_1 _2966_ (.CLK(net807),
    .D(net299),
    .Q(net561));
 sky130_fd_sc_hd__dfxtp_1 _2967_ (.CLK(net808),
    .D(net300),
    .Q(net468));
 sky130_fd_sc_hd__dfxtp_1 _2968_ (.CLK(net809),
    .D(net301),
    .Q(net469));
 sky130_fd_sc_hd__dfxtp_1 _2969_ (.CLK(net810),
    .D(net302),
    .Q(net470));
 sky130_fd_sc_hd__dfxtp_1 _2970_ (.CLK(net811),
    .D(net303),
    .Q(net471));
 sky130_fd_sc_hd__dfxtp_1 _2971_ (.CLK(net812),
    .D(net304),
    .Q(net472));
 sky130_fd_sc_hd__dfxtp_1 _2972_ (.CLK(net813),
    .D(net305),
    .Q(net473));
 sky130_fd_sc_hd__dfxtp_2 _2973_ (.CLK(net814),
    .D(net276),
    .Q(net474));
 sky130_fd_sc_hd__dfxtp_2 _2974_ (.CLK(net815),
    .D(net277),
    .Q(net475));
 sky130_fd_sc_hd__dfxtp_2 _2975_ (.CLK(net816),
    .D(net278),
    .Q(net476));
 sky130_fd_sc_hd__dfxtp_2 _2976_ (.CLK(net817),
    .D(net279),
    .Q(net477));
 sky130_fd_sc_hd__dfxtp_2 _2977_ (.CLK(net818),
    .D(net280),
    .Q(net479));
 sky130_fd_sc_hd__dfxtp_2 _2978_ (.CLK(net819),
    .D(net281),
    .Q(net480));
 sky130_fd_sc_hd__dfxtp_2 _2979_ (.CLK(net820),
    .D(net282),
    .Q(net481));
 sky130_fd_sc_hd__dfxtp_2 _2980_ (.CLK(net821),
    .D(net283),
    .Q(net482));
 sky130_fd_sc_hd__dfxtp_2 _2981_ (.CLK(net822),
    .D(net284),
    .Q(net483));
 sky130_fd_sc_hd__dfxtp_2 _2982_ (.CLK(net823),
    .D(net285),
    .Q(net484));
 sky130_fd_sc_hd__dfxtp_2 _2983_ (.CLK(net824),
    .D(net287),
    .Q(net485));
 sky130_fd_sc_hd__dfxtp_2 _2984_ (.CLK(net825),
    .D(net288),
    .Q(net486));
 sky130_fd_sc_hd__dfxtp_2 _2985_ (.CLK(net826),
    .D(net289),
    .Q(net487));
 sky130_fd_sc_hd__dfxtp_2 _2986_ (.CLK(net827),
    .D(net290),
    .Q(net488));
 sky130_fd_sc_hd__dfxtp_2 _2987_ (.CLK(net828),
    .D(net291),
    .Q(net490));
 sky130_fd_sc_hd__dfxtp_2 _2988_ (.CLK(net829),
    .D(net292),
    .Q(net491));
 sky130_fd_sc_hd__dfxtp_2 _2989_ (.CLK(net830),
    .D(net293),
    .Q(net492));
 sky130_fd_sc_hd__dfxtp_2 _2990_ (.CLK(net831),
    .D(net294),
    .Q(net493));
 sky130_fd_sc_hd__dfxtp_2 _2991_ (.CLK(net832),
    .D(net295),
    .Q(net494));
 sky130_fd_sc_hd__dfxtp_2 _2992_ (.CLK(net833),
    .D(net296),
    .Q(net495));
 sky130_fd_sc_hd__dfxtp_2 _2993_ (.CLK(net834),
    .D(net298),
    .Q(net496));
 sky130_fd_sc_hd__dfrtp_1 _2994_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0352_),
    .RESET_B(net600),
    .Q(net308));
 sky130_fd_sc_hd__dfrtp_1 _2995_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0353_),
    .RESET_B(net600),
    .Q(net319));
 sky130_fd_sc_hd__dfrtp_1 _2996_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0354_),
    .RESET_B(net600),
    .Q(net323));
 sky130_fd_sc_hd__dfrtp_1 _2997_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0355_),
    .RESET_B(net617),
    .Q(net324));
 sky130_fd_sc_hd__dfrtp_1 _2998_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0356_),
    .RESET_B(net617),
    .Q(net325));
 sky130_fd_sc_hd__dfrtp_1 _2999_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0357_),
    .RESET_B(net617),
    .Q(net326));
 sky130_fd_sc_hd__dfrtp_1 _3000_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0358_),
    .RESET_B(net617),
    .Q(net327));
 sky130_fd_sc_hd__dfrtp_1 _3001_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0359_),
    .RESET_B(net617),
    .Q(net328));
 sky130_fd_sc_hd__dfrtp_1 _3002_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0360_),
    .RESET_B(net617),
    .Q(net329));
 sky130_fd_sc_hd__dfrtp_1 _3003_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0361_),
    .RESET_B(net617),
    .Q(net330));
 sky130_fd_sc_hd__dfrtp_1 _3004_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0362_),
    .RESET_B(net617),
    .Q(net309));
 sky130_fd_sc_hd__dfrtp_1 _3005_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0363_),
    .RESET_B(net618),
    .Q(net310));
 sky130_fd_sc_hd__dfrtp_1 _3006_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0364_),
    .RESET_B(net620),
    .Q(net311));
 sky130_fd_sc_hd__dfrtp_1 _3007_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0365_),
    .RESET_B(net620),
    .Q(net312));
 sky130_fd_sc_hd__dfrtp_1 _3008_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0366_),
    .RESET_B(net620),
    .Q(net313));
 sky130_fd_sc_hd__dfrtp_1 _3009_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0367_),
    .RESET_B(net620),
    .Q(net314));
 sky130_fd_sc_hd__dfrtp_1 _3010_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0368_),
    .RESET_B(net620),
    .Q(net315));
 sky130_fd_sc_hd__dfrtp_1 _3011_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0369_),
    .RESET_B(net620),
    .Q(net316));
 sky130_fd_sc_hd__dfrtp_1 _3012_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0370_),
    .RESET_B(net622),
    .Q(net317));
 sky130_fd_sc_hd__dfrtp_1 _3013_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0371_),
    .RESET_B(net628),
    .Q(net318));
 sky130_fd_sc_hd__dfrtp_1 _3014_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0372_),
    .RESET_B(net628),
    .Q(net320));
 sky130_fd_sc_hd__dfrtp_1 _3015_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0373_),
    .RESET_B(net628),
    .Q(net321));
 sky130_fd_sc_hd__dfrtp_1 _3016_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0374_),
    .RESET_B(net628),
    .Q(net322));
 sky130_fd_sc_hd__dfrtp_2 _3017_ (.CLK(net835),
    .D(_0000_),
    .RESET_B(_0202_),
    .Q(prog_wea));
 sky130_fd_sc_hd__dfrtp_4 _3018_ (.CLK(net836),
    .D(_0375_),
    .RESET_B(_0204_),
    .Q(net563));
 sky130_fd_sc_hd__dfrtp_2 _3019_ (.CLK(net837),
    .D(_0376_),
    .RESET_B(_0206_),
    .Q(prog_h_addr0));
 sky130_fd_sc_hd__dfrtp_4 _3020_ (.CLK(net838),
    .D(_0377_),
    .RESET_B(_0208_),
    .Q(net383));
 sky130_fd_sc_hd__dfrtp_4 _3021_ (.CLK(net839),
    .D(_0378_),
    .RESET_B(_0210_),
    .Q(net384));
 sky130_fd_sc_hd__dfrtp_4 _3022_ (.CLK(net840),
    .D(_0379_),
    .RESET_B(_0212_),
    .Q(net385));
 sky130_fd_sc_hd__dfrtp_4 _3023_ (.CLK(net841),
    .D(_0380_),
    .RESET_B(_0214_),
    .Q(net386));
 sky130_fd_sc_hd__dfrtp_4 _3024_ (.CLK(net842),
    .D(_0381_),
    .RESET_B(_0216_),
    .Q(net387));
 sky130_fd_sc_hd__dfrtp_4 _3025_ (.CLK(net843),
    .D(_0382_),
    .RESET_B(_0218_),
    .Q(net388));
 sky130_fd_sc_hd__dfrtp_4 _3026_ (.CLK(net844),
    .D(_0383_),
    .RESET_B(_0220_),
    .Q(net389));
 sky130_fd_sc_hd__dfrtp_4 _3027_ (.CLK(net845),
    .D(_0384_),
    .RESET_B(_0222_),
    .Q(net390));
 sky130_fd_sc_hd__dfrtp_4 _3028_ (.CLK(net846),
    .D(_0385_),
    .RESET_B(_0224_),
    .Q(net392));
 sky130_fd_sc_hd__dfrtp_4 _3029_ (.CLK(net847),
    .D(_0386_),
    .RESET_B(_0226_),
    .Q(net403));
 sky130_fd_sc_hd__dfrtp_4 _3030_ (.CLK(net848),
    .D(_0387_),
    .RESET_B(_0228_),
    .Q(net414));
 sky130_fd_sc_hd__dfrtp_4 _3031_ (.CLK(net849),
    .D(_0388_),
    .RESET_B(_0230_),
    .Q(net417));
 sky130_fd_sc_hd__dfrtp_4 _3032_ (.CLK(net850),
    .D(_0389_),
    .RESET_B(_0232_),
    .Q(net418));
 sky130_fd_sc_hd__dfrtp_4 _3033_ (.CLK(net851),
    .D(_0390_),
    .RESET_B(_0234_),
    .Q(net419));
 sky130_fd_sc_hd__dfrtp_4 _3034_ (.CLK(net852),
    .D(_0391_),
    .RESET_B(_0236_),
    .Q(net420));
 sky130_fd_sc_hd__dfrtp_4 _3035_ (.CLK(net853),
    .D(_0392_),
    .RESET_B(_0238_),
    .Q(net421));
 sky130_fd_sc_hd__dfrtp_4 _3036_ (.CLK(net854),
    .D(_0393_),
    .RESET_B(_0240_),
    .Q(net422));
 sky130_fd_sc_hd__dfrtp_4 _3037_ (.CLK(net855),
    .D(_0394_),
    .RESET_B(_0242_),
    .Q(net423));
 sky130_fd_sc_hd__dfrtp_4 _3038_ (.CLK(net856),
    .D(_0395_),
    .RESET_B(_0244_),
    .Q(net393));
 sky130_fd_sc_hd__dfrtp_4 _3039_ (.CLK(net857),
    .D(_0396_),
    .RESET_B(_0246_),
    .Q(net394));
 sky130_fd_sc_hd__dfrtp_4 _3040_ (.CLK(net858),
    .D(_0397_),
    .RESET_B(_0248_),
    .Q(net395));
 sky130_fd_sc_hd__dfrtp_4 _3041_ (.CLK(net859),
    .D(_0398_),
    .RESET_B(_0250_),
    .Q(net396));
 sky130_fd_sc_hd__dfrtp_4 _3042_ (.CLK(net860),
    .D(_0399_),
    .RESET_B(_0252_),
    .Q(net397));
 sky130_fd_sc_hd__dfrtp_4 _3043_ (.CLK(net861),
    .D(_0400_),
    .RESET_B(_0254_),
    .Q(net398));
 sky130_fd_sc_hd__dfrtp_4 _3044_ (.CLK(net862),
    .D(_0401_),
    .RESET_B(_0256_),
    .Q(net399));
 sky130_fd_sc_hd__dfrtp_4 _3045_ (.CLK(net863),
    .D(_0402_),
    .RESET_B(_0258_),
    .Q(net400));
 sky130_fd_sc_hd__dfrtp_4 _3046_ (.CLK(net864),
    .D(_0403_),
    .RESET_B(_0260_),
    .Q(net401));
 sky130_fd_sc_hd__dfrtp_4 _3047_ (.CLK(net865),
    .D(_0404_),
    .RESET_B(_0262_),
    .Q(net402));
 sky130_fd_sc_hd__dfrtp_4 _3048_ (.CLK(net866),
    .D(_0405_),
    .RESET_B(_0264_),
    .Q(net404));
 sky130_fd_sc_hd__dfrtp_4 _3049_ (.CLK(net867),
    .D(_0406_),
    .RESET_B(_0266_),
    .Q(net405));
 sky130_fd_sc_hd__dfrtp_4 _3050_ (.CLK(net868),
    .D(_0407_),
    .RESET_B(_0268_),
    .Q(net406));
 sky130_fd_sc_hd__dfrtp_4 _3051_ (.CLK(net869),
    .D(_0408_),
    .RESET_B(_0270_),
    .Q(net407));
 sky130_fd_sc_hd__dfrtp_4 _3052_ (.CLK(net870),
    .D(_0409_),
    .RESET_B(_0272_),
    .Q(net408));
 sky130_fd_sc_hd__dfrtp_4 _3053_ (.CLK(net871),
    .D(_0410_),
    .RESET_B(_0274_),
    .Q(net409));
 sky130_fd_sc_hd__dfrtp_4 _3054_ (.CLK(net872),
    .D(_0411_),
    .RESET_B(_0276_),
    .Q(net410));
 sky130_fd_sc_hd__dfrtp_4 _3055_ (.CLK(net873),
    .D(_0412_),
    .RESET_B(_0278_),
    .Q(net411));
 sky130_fd_sc_hd__dfrtp_4 _3056_ (.CLK(net694),
    .D(_0413_),
    .RESET_B(_0280_),
    .Q(net412));
 sky130_fd_sc_hd__dfrtp_4 _3057_ (.CLK(net695),
    .D(_0414_),
    .RESET_B(_0282_),
    .Q(net413));
 sky130_fd_sc_hd__dfrtp_4 _3058_ (.CLK(net696),
    .D(_0415_),
    .RESET_B(_0284_),
    .Q(net415));
 sky130_fd_sc_hd__dfrtp_4 _3059_ (.CLK(net697),
    .D(_0416_),
    .RESET_B(_0286_),
    .Q(net416));
 sky130_fd_sc_hd__dfxtp_1 _3060_ (.CLK(net698),
    .D(net136),
    .Q(net467));
 sky130_fd_sc_hd__dfxtp_1 _3061_ (.CLK(net699),
    .D(net147),
    .Q(net505));
 sky130_fd_sc_hd__dfxtp_1 _3062_ (.CLK(net700),
    .D(net158),
    .Q(net516));
 sky130_fd_sc_hd__dfxtp_1 _3063_ (.CLK(net701),
    .D(net161),
    .Q(net527));
 sky130_fd_sc_hd__dfxtp_1 _3064_ (.CLK(net702),
    .D(net162),
    .Q(net538));
 sky130_fd_sc_hd__dfxtp_1 _3065_ (.CLK(net703),
    .D(net163),
    .Q(net549));
 sky130_fd_sc_hd__dfxtp_1 _3066_ (.CLK(net704),
    .D(net164),
    .Q(net554));
 sky130_fd_sc_hd__dfxtp_1 _3067_ (.CLK(net705),
    .D(net165),
    .Q(net555));
 sky130_fd_sc_hd__dfxtp_1 _3068_ (.CLK(net706),
    .D(net166),
    .Q(net556));
 sky130_fd_sc_hd__dfxtp_1 _3069_ (.CLK(net707),
    .D(net167),
    .Q(net562));
 sky130_fd_sc_hd__dfxtp_1 _3070_ (.CLK(net708),
    .D(net137),
    .Q(net478));
 sky130_fd_sc_hd__dfxtp_1 _3071_ (.CLK(net709),
    .D(net138),
    .Q(net489));
 sky130_fd_sc_hd__dfxtp_1 _3072_ (.CLK(net710),
    .D(net139),
    .Q(net497));
 sky130_fd_sc_hd__dfxtp_1 _3073_ (.CLK(net711),
    .D(net140),
    .Q(net498));
 sky130_fd_sc_hd__dfxtp_1 _3074_ (.CLK(net712),
    .D(net141),
    .Q(net499));
 sky130_fd_sc_hd__dfxtp_1 _3075_ (.CLK(net713),
    .D(net142),
    .Q(net500));
 sky130_fd_sc_hd__dfxtp_1 _3076_ (.CLK(net714),
    .D(net143),
    .Q(net501));
 sky130_fd_sc_hd__dfxtp_1 _3077_ (.CLK(net715),
    .D(net144),
    .Q(net502));
 sky130_fd_sc_hd__dfxtp_1 _3078_ (.CLK(net716),
    .D(net145),
    .Q(net503));
 sky130_fd_sc_hd__dfxtp_1 _3079_ (.CLK(net717),
    .D(net146),
    .Q(net504));
 sky130_fd_sc_hd__dfxtp_1 _3080_ (.CLK(net718),
    .D(net148),
    .Q(net506));
 sky130_fd_sc_hd__dfxtp_1 _3081_ (.CLK(net719),
    .D(net149),
    .Q(net507));
 sky130_fd_sc_hd__dfxtp_1 _3082_ (.CLK(net720),
    .D(net150),
    .Q(net508));
 sky130_fd_sc_hd__dfxtp_1 _3083_ (.CLK(net721),
    .D(net151),
    .Q(net509));
 sky130_fd_sc_hd__dfxtp_1 _3084_ (.CLK(net722),
    .D(net152),
    .Q(net510));
 sky130_fd_sc_hd__dfxtp_1 _3085_ (.CLK(net723),
    .D(net153),
    .Q(net511));
 sky130_fd_sc_hd__dfxtp_1 _3086_ (.CLK(net724),
    .D(net154),
    .Q(net512));
 sky130_fd_sc_hd__dfxtp_1 _3087_ (.CLK(net725),
    .D(net155),
    .Q(net513));
 sky130_fd_sc_hd__dfxtp_1 _3088_ (.CLK(net726),
    .D(net156),
    .Q(net514));
 sky130_fd_sc_hd__dfxtp_1 _3089_ (.CLK(net727),
    .D(net157),
    .Q(net515));
 sky130_fd_sc_hd__dfxtp_1 _3090_ (.CLK(net728),
    .D(net159),
    .Q(net517));
 sky130_fd_sc_hd__dfxtp_1 _3091_ (.CLK(net729),
    .D(net160),
    .Q(net518));
 sky130_fd_sc_hd__dfxtp_1 _3092_ (.CLK(net730),
    .D(net104),
    .Q(net519));
 sky130_fd_sc_hd__dfxtp_1 _3093_ (.CLK(net731),
    .D(net115),
    .Q(net520));
 sky130_fd_sc_hd__dfxtp_1 _3094_ (.CLK(net732),
    .D(net126),
    .Q(net521));
 sky130_fd_sc_hd__dfxtp_1 _3095_ (.CLK(net733),
    .D(net129),
    .Q(net522));
 sky130_fd_sc_hd__dfxtp_1 _3096_ (.CLK(net734),
    .D(net130),
    .Q(net523));
 sky130_fd_sc_hd__dfxtp_1 _3097_ (.CLK(net735),
    .D(net131),
    .Q(net524));
 sky130_fd_sc_hd__dfxtp_1 _3098_ (.CLK(net736),
    .D(net132),
    .Q(net525));
 sky130_fd_sc_hd__dfxtp_1 _3099_ (.CLK(net737),
    .D(net133),
    .Q(net526));
 sky130_fd_sc_hd__dfxtp_1 _3100_ (.CLK(net738),
    .D(net134),
    .Q(net528));
 sky130_fd_sc_hd__dfxtp_1 _3101_ (.CLK(net739),
    .D(net135),
    .Q(net529));
 sky130_fd_sc_hd__dfxtp_1 _3102_ (.CLK(net740),
    .D(net105),
    .Q(net530));
 sky130_fd_sc_hd__dfxtp_1 _3103_ (.CLK(net741),
    .D(net106),
    .Q(net531));
 sky130_fd_sc_hd__dfxtp_1 _3104_ (.CLK(net742),
    .D(net107),
    .Q(net532));
 sky130_fd_sc_hd__dfxtp_1 _3105_ (.CLK(net743),
    .D(net108),
    .Q(net533));
 sky130_fd_sc_hd__dfxtp_1 _3106_ (.CLK(net744),
    .D(net109),
    .Q(net534));
 sky130_fd_sc_hd__dfxtp_1 _3107_ (.CLK(net745),
    .D(net110),
    .Q(net535));
 sky130_fd_sc_hd__dfxtp_1 _3108_ (.CLK(net746),
    .D(net111),
    .Q(net536));
 sky130_fd_sc_hd__dfxtp_1 _3109_ (.CLK(net747),
    .D(net112),
    .Q(net537));
 sky130_fd_sc_hd__dfxtp_1 _3110_ (.CLK(net748),
    .D(net113),
    .Q(net539));
 sky130_fd_sc_hd__dfxtp_1 _3111_ (.CLK(net749),
    .D(net114),
    .Q(net540));
 sky130_fd_sc_hd__dfxtp_1 _3112_ (.CLK(net750),
    .D(net116),
    .Q(net541));
 sky130_fd_sc_hd__dfxtp_1 _3113_ (.CLK(net751),
    .D(net117),
    .Q(net542));
 sky130_fd_sc_hd__dfxtp_1 _3114_ (.CLK(net752),
    .D(net118),
    .Q(net543));
 sky130_fd_sc_hd__dfxtp_1 _3115_ (.CLK(net753),
    .D(net119),
    .Q(net544));
 sky130_fd_sc_hd__dfxtp_1 _3116_ (.CLK(net686),
    .D(net120),
    .Q(net545));
 sky130_fd_sc_hd__dfxtp_1 _3117_ (.CLK(net687),
    .D(net121),
    .Q(net546));
 sky130_fd_sc_hd__dfxtp_1 _3118_ (.CLK(net688),
    .D(net122),
    .Q(net547));
 sky130_fd_sc_hd__dfxtp_1 _3119_ (.CLK(net689),
    .D(net123),
    .Q(net548));
 sky130_fd_sc_hd__dfxtp_1 _3120_ (.CLK(net690),
    .D(net124),
    .Q(net550));
 sky130_fd_sc_hd__dfxtp_1 _3121_ (.CLK(net691),
    .D(net125),
    .Q(net551));
 sky130_fd_sc_hd__dfxtp_1 _3122_ (.CLK(net692),
    .D(net127),
    .Q(net552));
 sky130_fd_sc_hd__dfxtp_1 _3123_ (.CLK(net693),
    .D(net128),
    .Q(net553));
 sky130_fd_sc_hd__dfstp_1 _3124_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0016_),
    .SET_B(net621),
    .Q(\i_ca.ca_match_hs_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3125_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0004_),
    .RESET_B(net619),
    .Q(\i_ca.ca_match_hs_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3126_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0017_),
    .RESET_B(net619),
    .Q(\i_ca.ca_match_hs_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3127_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0417_),
    .RESET_B(net614),
    .Q(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3128_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0418_),
    .RESET_B(net614),
    .Q(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3129_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0419_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3130_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0420_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3131_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0421_),
    .RESET_B(net598),
    .Q(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3132_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0422_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3133_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0423_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3134_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0424_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_add_fill[8] ));
 sky130_fd_sc_hd__dfrtp_4 _3135_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0425_),
    .RESET_B(net623),
    .Q(\i_ca.ca_wr_add_start[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3136_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0426_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_add_start[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3137_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0427_),
    .RESET_B(net615),
    .Q(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3138_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0428_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_add_start[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3139_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0429_),
    .RESET_B(net623),
    .Q(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3140_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0430_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3141_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0431_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_add_start[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3142_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0432_),
    .RESET_B(net615),
    .Q(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__dfrtp_2 _3143_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0433_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_add_start[8] ));
 sky130_fd_sc_hd__dfstp_1 _3144_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0006_),
    .SET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3145_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0018_),
    .RESET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3146_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0019_),
    .RESET_B(net616),
    .Q(\i_ca.ca_rd_fsm_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3147_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0007_),
    .RESET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3148_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0020_),
    .RESET_B(net612),
    .Q(\i_ca.ca_rd_fsm_state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3149_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0021_),
    .RESET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3150_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0022_),
    .RESET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3151_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0008_),
    .RESET_B(net615),
    .Q(\i_ca.ca_rd_fsm_state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3152_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0009_),
    .RESET_B(net613),
    .Q(\i_ca.ca_rd_fsm_state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3153_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0434_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3154_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0435_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3155_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0436_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3156_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0437_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3157_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0438_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3158_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0439_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3159_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0440_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3160_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0441_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3161_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0442_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_dina[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3162_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0443_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3163_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0444_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3164_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0445_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3165_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0446_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3166_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0447_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[13] ));
 sky130_fd_sc_hd__dfrtp_1 _3167_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0448_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3168_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0449_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3169_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0450_),
    .RESET_B(net610),
    .Q(\i_ca.ca_wr_dina[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3170_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0451_),
    .RESET_B(net608),
    .Q(\i_ca.ca_wr_dina[17] ));
 sky130_fd_sc_hd__dfrtp_1 _3171_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0452_),
    .RESET_B(net608),
    .Q(\i_ca.ca_wr_dina[18] ));
 sky130_fd_sc_hd__dfrtp_1 _3172_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0453_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_dina[19] ));
 sky130_fd_sc_hd__dfrtp_1 _3173_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0454_),
    .RESET_B(net608),
    .Q(\i_ca.ca_wr_dina[20] ));
 sky130_fd_sc_hd__dfrtp_1 _3174_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0455_),
    .RESET_B(net608),
    .Q(\i_ca.ca_wr_dina[21] ));
 sky130_fd_sc_hd__dfrtp_1 _3175_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0456_),
    .RESET_B(net608),
    .Q(\i_ca.ca_wr_dina[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3176_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0457_),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_dina[32] ));
 sky130_fd_sc_hd__dfrtp_4 _3177_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0038_),
    .RESET_B(net600),
    .Q(\i_ca.ca_time_const[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3178_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0049_),
    .RESET_B(net599),
    .Q(\i_ca.ca_time_const[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3179_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0053_),
    .RESET_B(net599),
    .Q(\i_ca.ca_time_const[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3180_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0054_),
    .RESET_B(net599),
    .Q(\i_ca.ca_time_const[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3181_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0055_),
    .RESET_B(net600),
    .Q(\i_ca.ca_time_const[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3182_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0056_),
    .RESET_B(net619),
    .Q(\i_ca.ca_time_const[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3183_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0057_),
    .RESET_B(net617),
    .Q(\i_ca.ca_time_const[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3184_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0058_),
    .RESET_B(net617),
    .Q(\i_ca.ca_time_const[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3185_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0059_),
    .RESET_B(net619),
    .Q(\i_ca.ca_time_const[8] ));
 sky130_fd_sc_hd__dfrtp_4 _3186_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0060_),
    .RESET_B(net619),
    .Q(\i_ca.ca_time_const[9] ));
 sky130_fd_sc_hd__dfrtp_4 _3187_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0039_),
    .RESET_B(net619),
    .Q(\i_ca.ca_time_const[10] ));
 sky130_fd_sc_hd__dfrtp_4 _3188_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0040_),
    .RESET_B(net618),
    .Q(\i_ca.ca_time_const[11] ));
 sky130_fd_sc_hd__dfrtp_4 _3189_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0041_),
    .RESET_B(net620),
    .Q(\i_ca.ca_time_const[12] ));
 sky130_fd_sc_hd__dfrtp_4 _3190_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0042_),
    .RESET_B(net618),
    .Q(\i_ca.ca_time_const[13] ));
 sky130_fd_sc_hd__dfrtp_4 _3191_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0043_),
    .RESET_B(net620),
    .Q(\i_ca.ca_time_const[14] ));
 sky130_fd_sc_hd__dfrtp_4 _3192_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0044_),
    .RESET_B(net620),
    .Q(\i_ca.ca_time_const[15] ));
 sky130_fd_sc_hd__dfrtp_4 _3193_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0045_),
    .RESET_B(net622),
    .Q(\i_ca.ca_time_const[16] ));
 sky130_fd_sc_hd__dfrtp_4 _3194_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0046_),
    .RESET_B(net622),
    .Q(\i_ca.ca_time_const[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3195_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0047_),
    .RESET_B(net628),
    .Q(\i_ca.ca_time_const[18] ));
 sky130_fd_sc_hd__dfrtp_4 _3196_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0048_),
    .RESET_B(net628),
    .Q(\i_ca.ca_time_const[19] ));
 sky130_fd_sc_hd__dfrtp_4 _3197_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0050_),
    .RESET_B(net631),
    .Q(\i_ca.ca_time_const[20] ));
 sky130_fd_sc_hd__dfrtp_4 _3198_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0051_),
    .RESET_B(net631),
    .Q(\i_ca.ca_time_const[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3199_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0052_),
    .RESET_B(net631),
    .Q(\i_ca.ca_time_const[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3200_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0458_),
    .RESET_B(net600),
    .Q(\i_ca.hs_write_tid_wr0_const[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3201_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0459_),
    .RESET_B(net600),
    .Q(\i_ca.hs_write_tid_wr0_const[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3202_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0460_),
    .RESET_B(net599),
    .Q(\i_ca.hs_write_tid_wr0_const[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3203_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(\i_ca.hs_ready_meta ),
    .RESET_B(net618),
    .Q(net331));
 sky130_fd_sc_hd__dfrtp_4 _3204_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0461_),
    .RESET_B(net600),
    .Q(\i_ca.hs_write_dbus_wr_data_const[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3205_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0462_),
    .RESET_B(net600),
    .Q(\i_ca.hs_write_dbus_wr_data_const[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3206_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0463_),
    .RESET_B(net599),
    .Q(\i_ca.hs_write_dbus_wr_data_const[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3207_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0464_),
    .RESET_B(net599),
    .Q(\i_ca.hs_write_dbus_wr_data_const[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3208_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0465_),
    .RESET_B(net600),
    .Q(\i_ca.hs_write_dbus_wr_data_const[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3209_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0466_),
    .RESET_B(net604),
    .Q(\i_ca.hs_write_dbus_wr_data_const[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3210_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0467_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3211_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0468_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3212_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0469_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[8] ));
 sky130_fd_sc_hd__dfrtp_4 _3213_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0470_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[9] ));
 sky130_fd_sc_hd__dfrtp_4 _3214_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0471_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[10] ));
 sky130_fd_sc_hd__dfrtp_4 _3215_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0472_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[11] ));
 sky130_fd_sc_hd__dfrtp_4 _3216_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0473_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[12] ));
 sky130_fd_sc_hd__dfrtp_4 _3217_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0474_),
    .RESET_B(net596),
    .Q(\i_ca.hs_write_dbus_wr_data_const[13] ));
 sky130_fd_sc_hd__dfrtp_4 _3218_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0475_),
    .RESET_B(net603),
    .Q(\i_ca.hs_write_dbus_wr_data_const[14] ));
 sky130_fd_sc_hd__dfrtp_4 _3219_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0476_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[15] ));
 sky130_fd_sc_hd__dfrtp_4 _3220_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0477_),
    .RESET_B(net599),
    .Q(\i_ca.hs_write_dbus_wr_data_const[16] ));
 sky130_fd_sc_hd__dfrtp_4 _3221_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0478_),
    .RESET_B(net598),
    .Q(\i_ca.hs_write_dbus_wr_data_const[17] ));
 sky130_fd_sc_hd__dfrtp_4 _3222_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0479_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[18] ));
 sky130_fd_sc_hd__dfrtp_4 _3223_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0480_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[19] ));
 sky130_fd_sc_hd__dfrtp_4 _3224_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0481_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[20] ));
 sky130_fd_sc_hd__dfrtp_4 _3225_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0482_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3226_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0483_),
    .RESET_B(net619),
    .Q(\i_ca.hs_write_dbus_wr_data_const[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3227_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0484_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[23] ));
 sky130_fd_sc_hd__dfrtp_4 _3228_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0485_),
    .RESET_B(net619),
    .Q(\i_ca.hs_write_dbus_wr_data_const[24] ));
 sky130_fd_sc_hd__dfrtp_4 _3229_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0486_),
    .RESET_B(net613),
    .Q(\i_ca.hs_write_dbus_wr_data_const[25] ));
 sky130_fd_sc_hd__dfrtp_4 _3230_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0487_),
    .RESET_B(net612),
    .Q(\i_ca.hs_write_dbus_wr_data_const[26] ));
 sky130_fd_sc_hd__dfrtp_4 _3231_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0488_),
    .RESET_B(net613),
    .Q(\i_ca.hs_write_dbus_wr_data_const[27] ));
 sky130_fd_sc_hd__dfrtp_4 _3232_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0489_),
    .RESET_B(net614),
    .Q(\i_ca.hs_write_dbus_wr_data_const[28] ));
 sky130_fd_sc_hd__dfrtp_4 _3233_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0490_),
    .RESET_B(net619),
    .Q(\i_ca.hs_write_dbus_wr_data_const[29] ));
 sky130_fd_sc_hd__dfrtp_4 _3234_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0491_),
    .RESET_B(net613),
    .Q(\i_ca.hs_write_dbus_wr_data_const[30] ));
 sky130_fd_sc_hd__dfrtp_1 _3235_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0492_),
    .RESET_B(net613),
    .Q(\i_ca.hs_write_dbus_wr_data_const[31] ));
 sky130_fd_sc_hd__dfrtp_1 _3236_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0493_),
    .RESET_B(net599),
    .Q(net306));
 sky130_fd_sc_hd__dfrtp_4 _3237_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0037_),
    .RESET_B(net598),
    .Q(\i_ca.ca_wr_et_const ));
 sky130_fd_sc_hd__dfrtp_4 _3238_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0036_),
    .RESET_B(net598),
    .Q(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__dfrtp_2 _3239_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net37),
    .RESET_B(net601),
    .Q(\i_ca.ca_dbus_valid_meta ));
 sky130_fd_sc_hd__dfrtp_4 _3240_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0494_),
    .RESET_B(net612),
    .Q(\i_ca.ca_wr_sync_update_done ));
 sky130_fd_sc_hd__dfrtp_1 _3241_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0030_),
    .RESET_B(net603),
    .Q(\i_ca.ca_compare_check ));
 sky130_fd_sc_hd__dfrtp_1 _3242_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0029_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_equal_high ));
 sky130_fd_sc_hd__dfrtp_1 _3243_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0032_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_lesser_high ));
 sky130_fd_sc_hd__dfrtp_1 _3244_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0028_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_lesser_low ));
 sky130_fd_sc_hd__dfrtp_4 _3245_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0495_),
    .RESET_B(net614),
    .Q(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__dfrtp_1 _3246_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0496_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_time[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3247_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0497_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3248_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0498_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[2] ));
 sky130_fd_sc_hd__dfrtp_2 _3249_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0499_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3250_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0500_),
    .RESET_B(net608),
    .Q(\i_ca.ca_insert_time[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3251_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0501_),
    .RESET_B(net607),
    .Q(\i_ca.ca_insert_time[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3252_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0502_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3253_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0503_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3254_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0504_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3255_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0505_),
    .RESET_B(net608),
    .Q(\i_ca.ca_insert_time[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3256_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0506_),
    .RESET_B(net608),
    .Q(\i_ca.ca_insert_time[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3257_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0507_),
    .RESET_B(net608),
    .Q(\i_ca.ca_insert_time[11] ));
 sky130_fd_sc_hd__dfrtp_1 _3258_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0508_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[12] ));
 sky130_fd_sc_hd__dfrtp_2 _3259_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0509_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[13] ));
 sky130_fd_sc_hd__dfrtp_4 _3260_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0510_),
    .RESET_B(net605),
    .Q(\i_ca.ca_insert_time[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3261_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0511_),
    .RESET_B(net609),
    .Q(\i_ca.ca_insert_time[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3262_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0512_),
    .RESET_B(net609),
    .Q(\i_ca.ca_insert_time[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3263_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0513_),
    .RESET_B(net608),
    .Q(\i_ca.ca_insert_time[17] ));
 sky130_fd_sc_hd__dfrtp_2 _3264_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0514_),
    .RESET_B(net609),
    .Q(\i_ca.ca_insert_time[18] ));
 sky130_fd_sc_hd__dfrtp_2 _3265_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0515_),
    .RESET_B(net603),
    .Q(\i_ca.ca_insert_time[19] ));
 sky130_fd_sc_hd__dfrtp_2 _3266_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0516_),
    .RESET_B(net603),
    .Q(\i_ca.ca_insert_time[20] ));
 sky130_fd_sc_hd__dfrtp_2 _3267_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0517_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_time[21] ));
 sky130_fd_sc_hd__dfrtp_4 _3268_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0518_),
    .RESET_B(net604),
    .Q(\i_ca.ca_insert_time[22] ));
 sky130_fd_sc_hd__dfrtp_4 _3269_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0519_),
    .RESET_B(net597),
    .Q(\i_ca.ca_ready ));
 sky130_fd_sc_hd__dfrtp_4 _3270_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0520_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_dina[23] ));
 sky130_fd_sc_hd__dfrtp_4 _3271_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0521_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_dina[24] ));
 sky130_fd_sc_hd__dfrtp_4 _3272_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0522_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_dina[25] ));
 sky130_fd_sc_hd__dfrtp_4 _3273_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0523_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_dina[26] ));
 sky130_fd_sc_hd__dfrtp_4 _3274_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0524_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_dina[27] ));
 sky130_fd_sc_hd__dfrtp_4 _3275_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0525_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_dina[28] ));
 sky130_fd_sc_hd__dfrtp_4 _3276_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0526_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_dina[29] ));
 sky130_fd_sc_hd__dfrtp_4 _3277_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0527_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_dina[30] ));
 sky130_fd_sc_hd__dfrtp_1 _3278_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0528_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_dina[31] ));
 sky130_fd_sc_hd__dfrtp_1 _3279_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0529_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_add_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3280_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0530_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_add_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3281_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0531_),
    .RESET_B(net611),
    .Q(\i_ca.ca_wr_add_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3282_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0532_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_add_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3283_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0533_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_add_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3284_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0534_),
    .RESET_B(net624),
    .Q(\i_ca.ca_wr_add_ptr[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3285_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0535_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_add_ptr[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3286_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0536_),
    .RESET_B(net605),
    .Q(\i_ca.ca_wr_add_ptr[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3287_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0537_),
    .RESET_B(net606),
    .Q(\i_ca.ca_wr_add_ptr[8] ));
 sky130_fd_sc_hd__dfrtp_4 _3288_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0031_),
    .RESET_B(net625),
    .Q(\i_ca.ca_end_of_wr_list ));
 sky130_fd_sc_hd__dfrtp_4 _3289_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0538_),
    .RESET_B(net614),
    .Q(\i_ca.ca_wr_add_start_marker ));
 sky130_fd_sc_hd__dfrtp_4 _3290_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0539_),
    .RESET_B(net611),
    .Q(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3291_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0540_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__dfrtp_4 _3292_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0541_),
    .RESET_B(net611),
    .Q(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3293_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0542_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3294_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0543_),
    .RESET_B(net611),
    .Q(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__dfrtp_4 _3295_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0544_),
    .RESET_B(net625),
    .Q(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__dfrtp_4 _3296_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0545_),
    .RESET_B(net609),
    .Q(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3297_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0546_),
    .RESET_B(net606),
    .Q(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3298_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0547_),
    .RESET_B(net606),
    .Q(\i_ca.ca_wr_add[8] ));
 sky130_fd_sc_hd__dfrtp_4 _3299_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0548_),
    .RESET_B(net613),
    .Q(\i_ca.ca_wr_sync_update ));
 sky130_fd_sc_hd__dfrtp_1 _3300_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_1438_),
    .RESET_B(net607),
    .Q(\i_ca.ca_wr_wea ));
 sky130_fd_sc_hd__dfstp_1 _3301_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0002_),
    .SET_B(net601),
    .Q(\i_ca.hs_state_write_const[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3302_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0014_),
    .RESET_B(net599),
    .Q(\i_ca.hs_state_write_const[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3303_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0003_),
    .RESET_B(net601),
    .Q(\i_ca.hs_state_write_const[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3304_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0015_),
    .RESET_B(net599),
    .Q(\i_ca.hs_state_write_const[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net72),
    .Q(\i_ca.ca_rd_doutb[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net83),
    .Q(\i_ca.ca_rd_doutb[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3307_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net94),
    .Q(\i_ca.ca_rd_doutb[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3308_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net97),
    .Q(\i_ca.ca_rd_doutb[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3309_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net98),
    .Q(\i_ca.ca_rd_doutb[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3310_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net99),
    .Q(\i_ca.ca_rd_doutb[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3311_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net100),
    .Q(\i_ca.ca_rd_doutb[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3312_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net101),
    .Q(\i_ca.ca_rd_doutb[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3313_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net102),
    .Q(\i_ca.ca_rd_doutb[8] ));
 sky130_fd_sc_hd__dfxtp_2 _3314_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net103),
    .Q(\i_ca.ca_rd_doutb[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3315_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net73),
    .Q(\i_ca.ca_rd_doutb[10] ));
 sky130_fd_sc_hd__dfxtp_2 _3316_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net74),
    .Q(\i_ca.ca_rd_doutb[11] ));
 sky130_fd_sc_hd__dfxtp_4 _3317_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net75),
    .Q(\i_ca.ca_rd_doutb[12] ));
 sky130_fd_sc_hd__dfxtp_2 _3318_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net76),
    .Q(\i_ca.ca_rd_doutb[13] ));
 sky130_fd_sc_hd__dfxtp_2 _3319_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net77),
    .Q(\i_ca.ca_rd_doutb[14] ));
 sky130_fd_sc_hd__dfxtp_2 _3320_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net78),
    .Q(\i_ca.ca_rd_doutb[15] ));
 sky130_fd_sc_hd__dfxtp_2 _3321_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net79),
    .Q(\i_ca.ca_rd_doutb[16] ));
 sky130_fd_sc_hd__dfxtp_2 _3322_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net80),
    .Q(\i_ca.ca_rd_doutb[17] ));
 sky130_fd_sc_hd__dfxtp_2 _3323_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net81),
    .Q(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__dfxtp_2 _3324_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net82),
    .Q(\i_ca.ca_rd_doutb[19] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net84),
    .Q(\i_ca.ca_rd_doutb[20] ));
 sky130_fd_sc_hd__dfxtp_2 _3326_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net85),
    .Q(\i_ca.ca_rd_doutb[21] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net86),
    .Q(\i_ca.ca_rd_doutb[22] ));
 sky130_fd_sc_hd__dfxtp_2 _3328_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net87),
    .Q(\i_ca.ca_rd_doutb[23] ));
 sky130_fd_sc_hd__dfxtp_2 _3329_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net88),
    .Q(\i_ca.ca_rd_doutb[24] ));
 sky130_fd_sc_hd__dfxtp_2 _3330_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net89),
    .Q(\i_ca.ca_rd_doutb[25] ));
 sky130_fd_sc_hd__dfxtp_2 _3331_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net90),
    .Q(\i_ca.ca_rd_doutb[26] ));
 sky130_fd_sc_hd__dfxtp_2 _3332_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net91),
    .Q(\i_ca.ca_rd_doutb[27] ));
 sky130_fd_sc_hd__dfxtp_2 _3333_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net92),
    .Q(\i_ca.ca_rd_doutb[28] ));
 sky130_fd_sc_hd__dfxtp_2 _3334_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net93),
    .Q(\i_ca.ca_rd_doutb[29] ));
 sky130_fd_sc_hd__dfxtp_4 _3335_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net95),
    .Q(\i_ca.ca_rd_doutb[30] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net96),
    .Q(\i_ca.ca_rd_doutb[32] ));
 sky130_fd_sc_hd__dfrtp_1 _3337_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0061_),
    .RESET_B(net619),
    .Q(\i_ca.ca_time_diff[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3338_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0062_),
    .RESET_B(net621),
    .Q(\i_ca.ca_time_diff[13] ));
 sky130_fd_sc_hd__dfrtp_1 _3339_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0063_),
    .RESET_B(net621),
    .Q(\i_ca.ca_time_diff[14] ));
 sky130_fd_sc_hd__dfrtp_1 _3340_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0064_),
    .RESET_B(net621),
    .Q(\i_ca.ca_time_diff[15] ));
 sky130_fd_sc_hd__dfrtp_1 _3341_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0065_),
    .RESET_B(net621),
    .Q(\i_ca.ca_time_diff[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3342_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0066_),
    .RESET_B(net627),
    .Q(\i_ca.ca_time_diff[17] ));
 sky130_fd_sc_hd__dfrtp_1 _3343_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0067_),
    .RESET_B(net627),
    .Q(\i_ca.ca_time_diff[18] ));
 sky130_fd_sc_hd__dfrtp_1 _3344_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0068_),
    .RESET_B(net627),
    .Q(\i_ca.ca_time_diff[19] ));
 sky130_fd_sc_hd__dfrtp_1 _3345_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0069_),
    .RESET_B(net629),
    .Q(\i_ca.ca_time_diff[20] ));
 sky130_fd_sc_hd__dfrtp_1 _3346_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0070_),
    .RESET_B(net630),
    .Q(\i_ca.ca_time_diff[21] ));
 sky130_fd_sc_hd__dfrtp_1 _3347_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0071_),
    .RESET_B(net630),
    .Q(\i_ca.ca_time_diff[22] ));
 sky130_fd_sc_hd__dfrtp_1 _3348_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0033_),
    .RESET_B(net621),
    .Q(\i_ca.ca_match_check ));
 sky130_fd_sc_hd__dfrtp_1 _3349_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0034_),
    .RESET_B(net615),
    .Q(\i_ca.ca_match_req ));
 sky130_fd_sc_hd__dfrtp_4 _3350_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net876),
    .RESET_B(net630),
    .Q(\i_ca.ca_rd_doutb_32 ));
 sky130_fd_sc_hd__dfrtp_1 _3351_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0035_),
    .RESET_B(net612),
    .Q(\i_ca.ca_rd_doutb_31_23 ));
 sky130_fd_sc_hd__dfrtp_1 _3352_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0549_),
    .RESET_B(net624),
    .Q(\i_ca.ca_rd_add[0] ));
 sky130_fd_sc_hd__dfrtp_1 _3353_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0550_),
    .RESET_B(net625),
    .Q(\i_ca.ca_rd_add[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3354_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0551_),
    .RESET_B(net625),
    .Q(\i_ca.ca_rd_add[2] ));
 sky130_fd_sc_hd__dfrtp_1 _3355_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0552_),
    .RESET_B(net624),
    .Q(\i_ca.ca_rd_add[3] ));
 sky130_fd_sc_hd__dfrtp_1 _3356_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0553_),
    .RESET_B(net626),
    .Q(\i_ca.ca_rd_add[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3357_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0554_),
    .RESET_B(net624),
    .Q(\i_ca.ca_rd_add[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3358_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0555_),
    .RESET_B(net626),
    .Q(\i_ca.ca_rd_add[6] ));
 sky130_fd_sc_hd__dfrtp_1 _3359_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0556_),
    .RESET_B(net624),
    .Q(\i_ca.ca_rd_add[7] ));
 sky130_fd_sc_hd__dfrtp_4 _3360_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0557_),
    .RESET_B(net621),
    .Q(net307));
 sky130_fd_sc_hd__dfrtp_1 _3361_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0005_),
    .RESET_B(net615),
    .Q(\i_ca.ca_match_block_ack ));
 sky130_fd_sc_hd__dfrtp_2 _3362_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net38),
    .RESET_B(net620),
    .Q(\i_ca.ca_match_ack_meta ));
 sky130_fd_sc_hd__dfrtp_4 _3363_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0558_),
    .RESET_B(net616),
    .Q(net275));
 sky130_fd_sc_hd__dfrtp_4 _3364_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0559_),
    .RESET_B(net621),
    .Q(net286));
 sky130_fd_sc_hd__dfrtp_4 _3365_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0560_),
    .RESET_B(net626),
    .Q(net297));
 sky130_fd_sc_hd__dfrtp_4 _3366_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0561_),
    .RESET_B(net626),
    .Q(net299));
 sky130_fd_sc_hd__dfrtp_4 _3367_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0562_),
    .RESET_B(net626),
    .Q(net300));
 sky130_fd_sc_hd__dfrtp_4 _3368_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0563_),
    .RESET_B(net621),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_4 _3369_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0564_),
    .RESET_B(net627),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_4 _3370_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0565_),
    .RESET_B(net626),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_4 _3371_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0566_),
    .RESET_B(net627),
    .Q(net304));
 sky130_fd_sc_hd__dfrtp_4 _3372_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0567_),
    .RESET_B(net627),
    .Q(net305));
 sky130_fd_sc_hd__dfrtp_4 _3373_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0568_),
    .RESET_B(net627),
    .Q(net276));
 sky130_fd_sc_hd__dfrtp_4 _3374_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0569_),
    .RESET_B(net627),
    .Q(net277));
 sky130_fd_sc_hd__dfrtp_4 _3375_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0570_),
    .RESET_B(net627),
    .Q(net278));
 sky130_fd_sc_hd__dfrtp_4 _3376_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0571_),
    .RESET_B(net627),
    .Q(net279));
 sky130_fd_sc_hd__dfrtp_4 _3377_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0572_),
    .RESET_B(net628),
    .Q(net280));
 sky130_fd_sc_hd__dfrtp_4 _3378_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0573_),
    .RESET_B(net629),
    .Q(net281));
 sky130_fd_sc_hd__dfrtp_4 _3379_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0574_),
    .RESET_B(net628),
    .Q(net282));
 sky130_fd_sc_hd__dfrtp_4 _3380_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0575_),
    .RESET_B(net628),
    .Q(net283));
 sky130_fd_sc_hd__dfrtp_4 _3381_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0576_),
    .RESET_B(net629),
    .Q(net284));
 sky130_fd_sc_hd__dfrtp_4 _3382_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0577_),
    .RESET_B(net629),
    .Q(net285));
 sky130_fd_sc_hd__dfrtp_4 _3383_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0578_),
    .RESET_B(net630),
    .Q(net287));
 sky130_fd_sc_hd__dfrtp_4 _3384_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0579_),
    .RESET_B(net630),
    .Q(net288));
 sky130_fd_sc_hd__dfrtp_4 _3385_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0580_),
    .RESET_B(net630),
    .Q(net289));
 sky130_fd_sc_hd__dfrtp_4 _3386_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0581_),
    .RESET_B(net629),
    .Q(net290));
 sky130_fd_sc_hd__dfrtp_4 _3387_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0582_),
    .RESET_B(net629),
    .Q(net291));
 sky130_fd_sc_hd__dfrtp_4 _3388_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0583_),
    .RESET_B(net629),
    .Q(net292));
 sky130_fd_sc_hd__dfrtp_4 _3389_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0584_),
    .RESET_B(net629),
    .Q(net293));
 sky130_fd_sc_hd__dfrtp_4 _3390_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0585_),
    .RESET_B(net630),
    .Q(net294));
 sky130_fd_sc_hd__dfrtp_4 _3391_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0586_),
    .RESET_B(net629),
    .Q(net295));
 sky130_fd_sc_hd__dfrtp_4 _3392_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0587_),
    .RESET_B(net629),
    .Q(net296));
 sky130_fd_sc_hd__dfrtp_4 _3393_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0588_),
    .RESET_B(net621),
    .Q(net298));
 sky130_fd_sc_hd__dfxtp_2 _3394_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net40),
    .Q(\i_ca.ca_wr_douta[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3395_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net51),
    .Q(\i_ca.ca_wr_douta[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3396_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net62),
    .Q(\i_ca.ca_wr_douta[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3397_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net65),
    .Q(\i_ca.ca_wr_douta[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net66),
    .Q(\i_ca.ca_wr_douta[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net67),
    .Q(\i_ca.ca_wr_douta[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net68),
    .Q(\i_ca.ca_wr_douta[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net69),
    .Q(\i_ca.ca_wr_douta[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net70),
    .Q(\i_ca.ca_wr_douta[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net71),
    .Q(\i_ca.ca_wr_douta[9] ));
 sky130_fd_sc_hd__dfxtp_2 _3404_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net41),
    .Q(\i_ca.ca_wr_douta[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net42),
    .Q(\i_ca.ca_wr_douta[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net43),
    .Q(\i_ca.ca_wr_douta[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net44),
    .Q(\i_ca.ca_wr_douta[13] ));
 sky130_fd_sc_hd__dfxtp_2 _3408_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net45),
    .Q(\i_ca.ca_wr_douta[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net46),
    .Q(\i_ca.ca_wr_douta[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net47),
    .Q(\i_ca.ca_wr_douta[16] ));
 sky130_fd_sc_hd__dfxtp_1 _3411_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net48),
    .Q(\i_ca.ca_wr_douta[17] ));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net49),
    .Q(\i_ca.ca_wr_douta[18] ));
 sky130_fd_sc_hd__dfxtp_2 _3413_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net50),
    .Q(\i_ca.ca_wr_douta[19] ));
 sky130_fd_sc_hd__dfxtp_2 _3414_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net52),
    .Q(\i_ca.ca_wr_douta[20] ));
 sky130_fd_sc_hd__dfxtp_2 _3415_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net53),
    .Q(\i_ca.ca_wr_douta[21] ));
 sky130_fd_sc_hd__dfxtp_4 _3416_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net54),
    .Q(\i_ca.ca_wr_douta[22] ));
 sky130_fd_sc_hd__dfxtp_2 _3417_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net55),
    .Q(\i_ca.ca_wr_douta[23] ));
 sky130_fd_sc_hd__dfxtp_2 _3418_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net56),
    .Q(\i_ca.ca_wr_douta[24] ));
 sky130_fd_sc_hd__dfxtp_2 _3419_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net57),
    .Q(\i_ca.ca_wr_douta[25] ));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net58),
    .Q(\i_ca.ca_wr_douta[26] ));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net59),
    .Q(\i_ca.ca_wr_douta[27] ));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net60),
    .Q(\i_ca.ca_wr_douta[28] ));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net61),
    .Q(\i_ca.ca_wr_douta[29] ));
 sky130_fd_sc_hd__dfxtp_2 _3424_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net63),
    .Q(\i_ca.ca_wr_douta[30] ));
 sky130_fd_sc_hd__dfxtp_4 _3425_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net64),
    .Q(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__dfstp_1 _3426_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net39),
    .SET_B(net618),
    .Q(\i_ca.hs_ready_meta ));
 sky130_fd_sc_hd__dfstp_4 _3427_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0010_),
    .SET_B(net614),
    .Q(\i_ca.ca_wr_fsm_state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _3428_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net879),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_fsm_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _3429_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0011_),
    .RESET_B(net596),
    .Q(\i_ca.ca_wr_fsm_state[2] ));
 sky130_fd_sc_hd__dfrtp_4 _3430_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\i_ca.ca_wr_fsm_state[13] ),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_fsm_state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _3431_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0025_),
    .RESET_B(net616),
    .Q(\i_ca.ca_wr_fsm_state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _3432_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0012_),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_fsm_state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _3433_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net875),
    .RESET_B(net596),
    .Q(\i_ca.ca_wr_fsm_state[6] ));
 sky130_fd_sc_hd__dfrtp_4 _3434_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0026_),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_fsm_state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _3435_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(\i_ca.ca_wr_fsm_state[12] ),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_fsm_state[8] ));
 sky130_fd_sc_hd__dfrtp_1 _3436_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0027_),
    .RESET_B(net614),
    .Q(\i_ca.ca_wr_fsm_state[9] ));
 sky130_fd_sc_hd__dfrtp_1 _3437_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0013_),
    .RESET_B(net602),
    .Q(\i_ca.ca_wr_fsm_state[10] ));
 sky130_fd_sc_hd__dfrtp_1 _3438_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(\i_ca.ca_wr_fsm_state[3] ),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_fsm_state[11] ));
 sky130_fd_sc_hd__dfrtp_2 _3439_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0023_),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_fsm_state[12] ));
 sky130_fd_sc_hd__dfrtp_1 _3440_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net880),
    .RESET_B(net603),
    .Q(\i_ca.ca_wr_fsm_state[13] ));
 sky130_fd_sc_hd__dfrtp_4 _3441_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0024_),
    .RESET_B(net614),
    .Q(\i_ca.ca_wr_fsm_state[14] ));
 sky130_fd_sc_hd__dfrtp_4 _3442_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net877),
    .RESET_B(net602),
    .Q(\i_ca.ca_wr_fsm_state[15] ));
 sky130_fd_sc_hd__dfrtp_4 _3443_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0001_),
    .RESET_B(net604),
    .Q(\i_ca.ca_wr_fsm_state[16] ));
 sky130_fd_sc_hd__dfrtp_1 _3444_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net878),
    .RESET_B(net597),
    .Q(\i_ca.ca_wr_fsm_state[17] ));
 sky130_fd_sc_hd__conb_1 cawb_675 (.HI(net675));
 sky130_fd_sc_hd__conb_1 cawb_676 (.HI(net676));
 sky130_fd_sc_hd__conb_1 cawb_677 (.HI(net677));
 sky130_fd_sc_hd__conb_1 cawb_678 (.HI(net678));
 sky130_fd_sc_hd__conb_1 cawb_679 (.HI(net679));
 sky130_fd_sc_hd__conb_1 cawb_680 (.HI(net680));
 sky130_fd_sc_hd__conb_1 cawb_681 (.HI(net681));
 sky130_fd_sc_hd__conb_1 cawb_682 (.HI(net682));
 sky130_fd_sc_hd__conb_1 cawb_683 (.HI(net683));
 sky130_fd_sc_hd__conb_1 cawb_684 (.HI(net684));
 sky130_fd_sc_hd__conb_1 cawb_685 (.HI(net685));
 sky130_fd_sc_hd__inv_2 _2325__1 (.A(clknet_1_1__leaf__0984_),
    .Y(net686));
 sky130_fd_sc_hd__conb_1 cawb_634 (.LO(net634));
 sky130_fd_sc_hd__conb_1 cawb_635 (.LO(net635));
 sky130_fd_sc_hd__conb_1 cawb_636 (.LO(net636));
 sky130_fd_sc_hd__conb_1 cawb_637 (.LO(net637));
 sky130_fd_sc_hd__conb_1 cawb_638 (.LO(net638));
 sky130_fd_sc_hd__conb_1 cawb_639 (.LO(net639));
 sky130_fd_sc_hd__conb_1 cawb_640 (.LO(net640));
 sky130_fd_sc_hd__conb_1 cawb_641 (.LO(net641));
 sky130_fd_sc_hd__conb_1 cawb_642 (.LO(net642));
 sky130_fd_sc_hd__conb_1 cawb_643 (.LO(net643));
 sky130_fd_sc_hd__conb_1 cawb_644 (.LO(net644));
 sky130_fd_sc_hd__conb_1 cawb_645 (.LO(net645));
 sky130_fd_sc_hd__conb_1 cawb_646 (.LO(net646));
 sky130_fd_sc_hd__conb_1 cawb_647 (.LO(net647));
 sky130_fd_sc_hd__conb_1 cawb_648 (.LO(net648));
 sky130_fd_sc_hd__conb_1 cawb_649 (.LO(net649));
 sky130_fd_sc_hd__conb_1 cawb_650 (.LO(net650));
 sky130_fd_sc_hd__conb_1 cawb_651 (.LO(net651));
 sky130_fd_sc_hd__conb_1 cawb_652 (.LO(net652));
 sky130_fd_sc_hd__conb_1 cawb_653 (.LO(net653));
 sky130_fd_sc_hd__conb_1 cawb_654 (.LO(net654));
 sky130_fd_sc_hd__conb_1 cawb_655 (.LO(net655));
 sky130_fd_sc_hd__conb_1 cawb_656 (.LO(net656));
 sky130_fd_sc_hd__conb_1 cawb_657 (.LO(net657));
 sky130_fd_sc_hd__conb_1 cawb_658 (.LO(net658));
 sky130_fd_sc_hd__conb_1 cawb_659 (.LO(net659));
 sky130_fd_sc_hd__conb_1 cawb_660 (.LO(net660));
 sky130_fd_sc_hd__conb_1 cawb_661 (.LO(net661));
 sky130_fd_sc_hd__conb_1 cawb_662 (.LO(net662));
 sky130_fd_sc_hd__conb_1 cawb_663 (.LO(net663));
 sky130_fd_sc_hd__conb_1 cawb_664 (.LO(net664));
 sky130_fd_sc_hd__conb_1 cawb_665 (.LO(net665));
 sky130_fd_sc_hd__conb_1 cawb_666 (.LO(net666));
 sky130_fd_sc_hd__conb_1 cawb_667 (.LO(net667));
 sky130_fd_sc_hd__conb_1 cawb_668 (.LO(net668));
 sky130_fd_sc_hd__conb_1 cawb_669 (.LO(net669));
 sky130_fd_sc_hd__conb_1 cawb_670 (.LO(net670));
 sky130_fd_sc_hd__conb_1 cawb_671 (.LO(net671));
 sky130_fd_sc_hd__conb_1 cawb_672 (.LO(net672));
 sky130_fd_sc_hd__conb_1 cawb_673 (.LO(net673));
 sky130_fd_sc_hd__conb_1 cawb_674 (.HI(net674));
 sky130_fd_sc_hd__buf_2 _3498_ (.A(clknet_opt_4_1_wb_clk_i),
    .X(net348));
 sky130_fd_sc_hd__buf_2 _3499_ (.A(clknet_leaf_26_wb_clk_i),
    .X(net349));
 sky130_fd_sc_hd__buf_2 _3500_ (.A(clknet_opt_3_2_wb_clk_i),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(net383),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 _3502_ (.A(net384),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 _3503_ (.A(net385),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 _3504_ (.A(net386),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(net387),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 _3506_ (.A(net388),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 _3507_ (.A(net389),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(net390),
    .X(net432));
 sky130_fd_sc_hd__buf_2 _3509_ (.A(clknet_opt_2_3_wb_clk_i),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(net392),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 _3511_ (.A(net403),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 _3512_ (.A(net414),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 _3513_ (.A(net417),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 _3514_ (.A(net418),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 _3515_ (.A(net419),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 _3516_ (.A(net420),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(net421),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 _3518_ (.A(net422),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(net423),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 _3520_ (.A(net393),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 _3521_ (.A(net394),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 _3522_ (.A(net395),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 _3523_ (.A(net396),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(net397),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 _3525_ (.A(net398),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 _3526_ (.A(net399),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 _3527_ (.A(net400),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 _3528_ (.A(net401),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 _3529_ (.A(net402),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 _3530_ (.A(net404),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 _3531_ (.A(net405),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 _3532_ (.A(net406),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 _3533_ (.A(net407),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 _3534_ (.A(net408),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 _3535_ (.A(net409),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 _3536_ (.A(net410),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 _3537_ (.A(net411),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 _3538_ (.A(net412),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 _3539_ (.A(net413),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 _3540_ (.A(net415),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_2 _3541_ (.A(net416),
    .X(net458));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ca_dbus_com),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ca_dbus_data[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(ca_dbus_data[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(ca_dbus_data[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(ca_dbus_data[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(ca_dbus_data[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ca_dbus_data[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ca_dbus_data[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ca_dbus_data[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(ca_dbus_data[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(ca_dbus_data[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(ca_dbus_data[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(ca_dbus_data[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(ca_dbus_data[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(ca_dbus_data[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(ca_dbus_data[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(ca_dbus_data[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(ca_dbus_data[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(ca_dbus_data[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(ca_dbus_data[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(ca_dbus_data[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(ca_dbus_data[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(ca_dbus_data[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(ca_dbus_data[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(ca_dbus_data[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(ca_dbus_data[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(ca_dbus_data[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(ca_dbus_data[4]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(ca_dbus_data[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(ca_dbus_data[6]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(ca_dbus_data[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(ca_dbus_data[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(ca_dbus_data[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(ca_dbus_tid[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(ca_dbus_tid[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(ca_dbus_tid[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(ca_dbus_valid),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(ca_match_ack),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(ca_time_ack),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(cubev_ca_dout0[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(cubev_ca_dout0[10]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(cubev_ca_dout0[11]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(cubev_ca_dout0[12]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(cubev_ca_dout0[13]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(cubev_ca_dout0[14]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(cubev_ca_dout0[15]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(cubev_ca_dout0[16]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(cubev_ca_dout0[17]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(cubev_ca_dout0[18]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(cubev_ca_dout0[19]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(cubev_ca_dout0[1]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(cubev_ca_dout0[20]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(cubev_ca_dout0[21]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(cubev_ca_dout0[22]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(cubev_ca_dout0[23]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(cubev_ca_dout0[24]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(cubev_ca_dout0[25]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(cubev_ca_dout0[26]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(cubev_ca_dout0[27]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(cubev_ca_dout0[28]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(cubev_ca_dout0[29]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(cubev_ca_dout0[2]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(cubev_ca_dout0[30]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(cubev_ca_dout0[31]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(cubev_ca_dout0[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(cubev_ca_dout0[4]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(cubev_ca_dout0[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(cubev_ca_dout0[6]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(cubev_ca_dout0[7]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(cubev_ca_dout0[8]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(cubev_ca_dout0[9]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(cubev_ca_dout1[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(cubev_ca_dout1[10]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(cubev_ca_dout1[11]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(cubev_ca_dout1[12]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(cubev_ca_dout1[13]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(cubev_ca_dout1[14]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(cubev_ca_dout1[15]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(cubev_ca_dout1[16]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(cubev_ca_dout1[17]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(cubev_ca_dout1[18]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(cubev_ca_dout1[19]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(cubev_ca_dout1[1]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(cubev_ca_dout1[20]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(cubev_ca_dout1[21]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(cubev_ca_dout1[22]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(cubev_ca_dout1[23]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(cubev_ca_dout1[24]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(cubev_ca_dout1[25]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(cubev_ca_dout1[26]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(cubev_ca_dout1[27]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(cubev_ca_dout1[28]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(cubev_ca_dout1[29]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(cubev_ca_dout1[2]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(cubev_ca_dout1[30]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(cubev_ca_dout1[31]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(cubev_ca_dout1[3]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(cubev_ca_dout1[4]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(cubev_ca_dout1[5]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(cubev_ca_dout1[6]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(cubev_ca_dout1[7]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(cubev_ca_dout1[8]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(cubev_ca_dout1[9]),
    .X(net103));
 sky130_fd_sc_hd__buf_6 input104 (.A(cubev_phi_dout0[0]),
    .X(net104));
 sky130_fd_sc_hd__buf_6 input105 (.A(cubev_phi_dout0[10]),
    .X(net105));
 sky130_fd_sc_hd__buf_6 input106 (.A(cubev_phi_dout0[11]),
    .X(net106));
 sky130_fd_sc_hd__buf_6 input107 (.A(cubev_phi_dout0[12]),
    .X(net107));
 sky130_fd_sc_hd__buf_6 input108 (.A(cubev_phi_dout0[13]),
    .X(net108));
 sky130_fd_sc_hd__buf_6 input109 (.A(cubev_phi_dout0[14]),
    .X(net109));
 sky130_fd_sc_hd__buf_6 input110 (.A(cubev_phi_dout0[15]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 input111 (.A(cubev_phi_dout0[16]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 input112 (.A(cubev_phi_dout0[17]),
    .X(net112));
 sky130_fd_sc_hd__buf_6 input113 (.A(cubev_phi_dout0[18]),
    .X(net113));
 sky130_fd_sc_hd__buf_6 input114 (.A(cubev_phi_dout0[19]),
    .X(net114));
 sky130_fd_sc_hd__buf_6 input115 (.A(cubev_phi_dout0[1]),
    .X(net115));
 sky130_fd_sc_hd__buf_6 input116 (.A(cubev_phi_dout0[20]),
    .X(net116));
 sky130_fd_sc_hd__buf_6 input117 (.A(cubev_phi_dout0[21]),
    .X(net117));
 sky130_fd_sc_hd__buf_6 input118 (.A(cubev_phi_dout0[22]),
    .X(net118));
 sky130_fd_sc_hd__buf_6 input119 (.A(cubev_phi_dout0[23]),
    .X(net119));
 sky130_fd_sc_hd__buf_6 input120 (.A(cubev_phi_dout0[24]),
    .X(net120));
 sky130_fd_sc_hd__buf_6 input121 (.A(cubev_phi_dout0[25]),
    .X(net121));
 sky130_fd_sc_hd__buf_6 input122 (.A(cubev_phi_dout0[26]),
    .X(net122));
 sky130_fd_sc_hd__buf_6 input123 (.A(cubev_phi_dout0[27]),
    .X(net123));
 sky130_fd_sc_hd__buf_6 input124 (.A(cubev_phi_dout0[28]),
    .X(net124));
 sky130_fd_sc_hd__buf_6 input125 (.A(cubev_phi_dout0[29]),
    .X(net125));
 sky130_fd_sc_hd__buf_6 input126 (.A(cubev_phi_dout0[2]),
    .X(net126));
 sky130_fd_sc_hd__buf_6 input127 (.A(cubev_phi_dout0[30]),
    .X(net127));
 sky130_fd_sc_hd__buf_6 input128 (.A(cubev_phi_dout0[31]),
    .X(net128));
 sky130_fd_sc_hd__buf_6 input129 (.A(cubev_phi_dout0[3]),
    .X(net129));
 sky130_fd_sc_hd__buf_6 input130 (.A(cubev_phi_dout0[4]),
    .X(net130));
 sky130_fd_sc_hd__buf_6 input131 (.A(cubev_phi_dout0[5]),
    .X(net131));
 sky130_fd_sc_hd__buf_6 input132 (.A(cubev_phi_dout0[6]),
    .X(net132));
 sky130_fd_sc_hd__buf_6 input133 (.A(cubev_phi_dout0[7]),
    .X(net133));
 sky130_fd_sc_hd__buf_6 input134 (.A(cubev_phi_dout0[8]),
    .X(net134));
 sky130_fd_sc_hd__buf_6 input135 (.A(cubev_phi_dout0[9]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(cubev_pli_dout0[0]),
    .X(net136));
 sky130_fd_sc_hd__buf_4 input137 (.A(cubev_pli_dout0[10]),
    .X(net137));
 sky130_fd_sc_hd__buf_4 input138 (.A(cubev_pli_dout0[11]),
    .X(net138));
 sky130_fd_sc_hd__buf_4 input139 (.A(cubev_pli_dout0[12]),
    .X(net139));
 sky130_fd_sc_hd__buf_4 input140 (.A(cubev_pli_dout0[13]),
    .X(net140));
 sky130_fd_sc_hd__buf_4 input141 (.A(cubev_pli_dout0[14]),
    .X(net141));
 sky130_fd_sc_hd__buf_4 input142 (.A(cubev_pli_dout0[15]),
    .X(net142));
 sky130_fd_sc_hd__buf_4 input143 (.A(cubev_pli_dout0[16]),
    .X(net143));
 sky130_fd_sc_hd__buf_4 input144 (.A(cubev_pli_dout0[17]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 input145 (.A(cubev_pli_dout0[18]),
    .X(net145));
 sky130_fd_sc_hd__buf_6 input146 (.A(cubev_pli_dout0[19]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(cubev_pli_dout0[1]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_8 input148 (.A(cubev_pli_dout0[20]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_8 input149 (.A(cubev_pli_dout0[21]),
    .X(net149));
 sky130_fd_sc_hd__buf_6 input150 (.A(cubev_pli_dout0[22]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_8 input151 (.A(cubev_pli_dout0[23]),
    .X(net151));
 sky130_fd_sc_hd__buf_6 input152 (.A(cubev_pli_dout0[24]),
    .X(net152));
 sky130_fd_sc_hd__buf_6 input153 (.A(cubev_pli_dout0[25]),
    .X(net153));
 sky130_fd_sc_hd__buf_6 input154 (.A(cubev_pli_dout0[26]),
    .X(net154));
 sky130_fd_sc_hd__buf_6 input155 (.A(cubev_pli_dout0[27]),
    .X(net155));
 sky130_fd_sc_hd__buf_6 input156 (.A(cubev_pli_dout0[28]),
    .X(net156));
 sky130_fd_sc_hd__buf_6 input157 (.A(cubev_pli_dout0[29]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(cubev_pli_dout0[2]),
    .X(net158));
 sky130_fd_sc_hd__buf_6 input159 (.A(cubev_pli_dout0[30]),
    .X(net159));
 sky130_fd_sc_hd__buf_6 input160 (.A(cubev_pli_dout0[31]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(cubev_pli_dout0[3]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(cubev_pli_dout0[4]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(cubev_pli_dout0[5]),
    .X(net163));
 sky130_fd_sc_hd__buf_4 input164 (.A(cubev_pli_dout0[6]),
    .X(net164));
 sky130_fd_sc_hd__buf_4 input165 (.A(cubev_pli_dout0[7]),
    .X(net165));
 sky130_fd_sc_hd__buf_4 input166 (.A(cubev_pli_dout0[8]),
    .X(net166));
 sky130_fd_sc_hd__buf_4 input167 (.A(cubev_pli_dout0[9]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(la_data_in[0]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(la_data_in[10]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(la_data_in[11]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(la_data_in[12]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 input172 (.A(la_data_in[13]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(la_data_in[14]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(la_data_in[15]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(la_data_in[16]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(la_data_in[17]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(la_data_in[18]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(la_data_in[19]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(la_data_in[1]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(la_data_in[20]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 input181 (.A(la_data_in[21]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(la_data_in[22]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(la_data_in[23]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(la_data_in[24]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(la_data_in[25]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(la_data_in[26]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(la_data_in[27]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(la_data_in[28]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(la_data_in[29]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(la_data_in[2]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(la_data_in[30]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(la_data_in[31]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 input193 (.A(la_data_in[32]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(la_data_in[33]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(la_data_in[34]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(la_data_in[35]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 input197 (.A(la_data_in[36]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(la_data_in[37]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(la_data_in[38]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(la_data_in[39]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(la_data_in[3]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(la_data_in[40]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(la_data_in[4]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(la_data_in[5]),
    .X(net204));
 sky130_fd_sc_hd__buf_4 input205 (.A(la_data_in[64]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(la_data_in[65]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 input207 (.A(la_data_in[6]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(la_data_in[7]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(la_data_in[8]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 input210 (.A(la_data_in[9]),
    .X(net210));
 sky130_fd_sc_hd__buf_6 input211 (.A(wb_rst_i),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 input212 (.A(wbs_adr_i[0]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(wbs_adr_i[10]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(wbs_adr_i[11]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(wbs_adr_i[16]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(wbs_adr_i[17]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(wbs_adr_i[18]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(wbs_adr_i[19]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(wbs_adr_i[1]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 input220 (.A(wbs_adr_i[20]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(wbs_adr_i[21]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(wbs_adr_i[22]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(wbs_adr_i[23]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(wbs_adr_i[24]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(wbs_adr_i[25]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(wbs_adr_i[26]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(wbs_adr_i[27]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(wbs_adr_i[28]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(wbs_adr_i[29]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(wbs_adr_i[2]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(wbs_adr_i[30]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(wbs_adr_i[31]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(wbs_adr_i[3]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(wbs_adr_i[4]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(wbs_adr_i[5]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(wbs_adr_i[6]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(wbs_adr_i[7]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(wbs_adr_i[8]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(wbs_adr_i[9]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(wbs_cyc_i),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(wbs_dat_i[0]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(wbs_dat_i[10]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(wbs_dat_i[11]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(wbs_dat_i[12]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 input245 (.A(wbs_dat_i[13]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(wbs_dat_i[14]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 input247 (.A(wbs_dat_i[15]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(wbs_dat_i[16]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(wbs_dat_i[17]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(wbs_dat_i[18]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(wbs_dat_i[19]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(wbs_dat_i[1]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(wbs_dat_i[20]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(wbs_dat_i[21]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(wbs_dat_i[22]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(wbs_dat_i[23]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 input257 (.A(wbs_dat_i[24]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(wbs_dat_i[25]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(wbs_dat_i[26]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 input260 (.A(wbs_dat_i[27]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 input261 (.A(wbs_dat_i[28]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input262 (.A(wbs_dat_i[29]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 input263 (.A(wbs_dat_i[2]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 input264 (.A(wbs_dat_i[30]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 input265 (.A(wbs_dat_i[31]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(wbs_dat_i[3]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 input267 (.A(wbs_dat_i[4]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 input268 (.A(wbs_dat_i[5]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(wbs_dat_i[6]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 input270 (.A(wbs_dat_i[7]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 input271 (.A(wbs_dat_i[8]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 input272 (.A(wbs_dat_i[9]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 input273 (.A(wbs_stb_i),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 input274 (.A(wbs_we_i),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(ca_command[0]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(ca_command[10]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .X(ca_command[11]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(ca_command[12]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .X(ca_command[13]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(ca_command[14]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(ca_command[15]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .X(ca_command[16]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(ca_command[17]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(ca_command[18]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(ca_command[19]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .X(ca_command[1]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .X(ca_command[20]));
 sky130_fd_sc_hd__clkbuf_4 output288 (.A(net288),
    .X(ca_command[21]));
 sky130_fd_sc_hd__clkbuf_4 output289 (.A(net289),
    .X(ca_command[22]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .X(ca_command[23]));
 sky130_fd_sc_hd__clkbuf_4 output291 (.A(net291),
    .X(ca_command[24]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .X(ca_command[25]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .X(ca_command[26]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .X(ca_command[27]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .X(ca_command[28]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .X(ca_command[29]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .X(ca_command[2]));
 sky130_fd_sc_hd__clkbuf_4 output298 (.A(net298),
    .X(ca_command[30]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .X(ca_command[3]));
 sky130_fd_sc_hd__clkbuf_4 output300 (.A(net300),
    .X(ca_command[4]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .X(ca_command[5]));
 sky130_fd_sc_hd__clkbuf_4 output302 (.A(net302),
    .X(ca_command[6]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .X(ca_command[7]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .X(ca_command[8]));
 sky130_fd_sc_hd__clkbuf_4 output305 (.A(net305),
    .X(ca_command[9]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .X(ca_dbus_ack));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .X(ca_match_valid));
 sky130_fd_sc_hd__clkbuf_4 output308 (.A(net308),
    .X(ca_time_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .X(ca_time_data[10]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .X(ca_time_data[11]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .X(ca_time_data[12]));
 sky130_fd_sc_hd__clkbuf_4 output312 (.A(net312),
    .X(ca_time_data[13]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .X(ca_time_data[14]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .X(ca_time_data[15]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .X(ca_time_data[16]));
 sky130_fd_sc_hd__clkbuf_4 output316 (.A(net316),
    .X(ca_time_data[17]));
 sky130_fd_sc_hd__clkbuf_4 output317 (.A(net317),
    .X(ca_time_data[18]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .X(ca_time_data[19]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .X(ca_time_data[1]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .X(ca_time_data[20]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .X(ca_time_data[21]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .X(ca_time_data[22]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .X(ca_time_data[2]));
 sky130_fd_sc_hd__clkbuf_4 output324 (.A(net324),
    .X(ca_time_data[3]));
 sky130_fd_sc_hd__clkbuf_4 output325 (.A(net325),
    .X(ca_time_data[4]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .X(ca_time_data[5]));
 sky130_fd_sc_hd__clkbuf_4 output327 (.A(net327),
    .X(ca_time_data[6]));
 sky130_fd_sc_hd__clkbuf_4 output328 (.A(net328),
    .X(ca_time_data[7]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .X(ca_time_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .X(ca_time_data[9]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .X(ca_time_valid));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .X(cubev_ca_addr0[0]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .X(cubev_ca_addr0[1]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .X(cubev_ca_addr0[2]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .X(cubev_ca_addr0[3]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .X(cubev_ca_addr0[4]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .X(cubev_ca_addr0[5]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .X(cubev_ca_addr0[6]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .X(cubev_ca_addr0[7]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .X(cubev_ca_addr1[0]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .X(cubev_ca_addr1[1]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .X(cubev_ca_addr1[2]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .X(cubev_ca_addr1[3]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .X(cubev_ca_addr1[4]));
 sky130_fd_sc_hd__clkbuf_4 output345 (.A(net345),
    .X(cubev_ca_addr1[5]));
 sky130_fd_sc_hd__clkbuf_4 output346 (.A(net346),
    .X(cubev_ca_addr1[6]));
 sky130_fd_sc_hd__clkbuf_4 output347 (.A(net347),
    .X(cubev_ca_addr1[7]));
 sky130_fd_sc_hd__clkbuf_1 output348 (.A(net348),
    .X(cubev_ca_clk0));
 sky130_fd_sc_hd__clkbuf_1 output349 (.A(net349),
    .X(cubev_ca_clk1));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .X(cubev_ca_din0[0]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .X(cubev_ca_din0[10]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .X(cubev_ca_din0[11]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .X(cubev_ca_din0[12]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .X(cubev_ca_din0[13]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .X(cubev_ca_din0[14]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(cubev_ca_din0[15]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .X(cubev_ca_din0[16]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .X(cubev_ca_din0[17]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .X(cubev_ca_din0[18]));
 sky130_fd_sc_hd__clkbuf_4 output360 (.A(net360),
    .X(cubev_ca_din0[19]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .X(cubev_ca_din0[1]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .X(cubev_ca_din0[20]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .X(cubev_ca_din0[21]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .X(cubev_ca_din0[22]));
 sky130_fd_sc_hd__clkbuf_4 output365 (.A(net365),
    .X(cubev_ca_din0[23]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .X(cubev_ca_din0[24]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .X(cubev_ca_din0[25]));
 sky130_fd_sc_hd__clkbuf_4 output368 (.A(net368),
    .X(cubev_ca_din0[26]));
 sky130_fd_sc_hd__clkbuf_4 output369 (.A(net369),
    .X(cubev_ca_din0[27]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .X(cubev_ca_din0[28]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .X(cubev_ca_din0[29]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .X(cubev_ca_din0[2]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .X(cubev_ca_din0[30]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .X(cubev_ca_din0[31]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .X(cubev_ca_din0[3]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .X(cubev_ca_din0[4]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .X(cubev_ca_din0[5]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .X(cubev_ca_din0[6]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .X(cubev_ca_din0[7]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .X(cubev_ca_din0[8]));
 sky130_fd_sc_hd__clkbuf_4 output381 (.A(net381),
    .X(cubev_ca_din0[9]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .X(cubev_ca_web0));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(cubev_phi_addr0[0]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(cubev_phi_addr0[1]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .X(cubev_phi_addr0[2]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .X(cubev_phi_addr0[3]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(cubev_phi_addr0[4]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .X(cubev_phi_addr0[5]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .X(cubev_phi_addr0[6]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .X(cubev_phi_addr0[7]));
 sky130_fd_sc_hd__clkbuf_1 output391 (.A(net391),
    .X(cubev_phi_clk0));
 sky130_fd_sc_hd__clkbuf_4 output392 (.A(net392),
    .X(cubev_phi_din0[0]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .X(cubev_phi_din0[10]));
 sky130_fd_sc_hd__clkbuf_4 output394 (.A(net394),
    .X(cubev_phi_din0[11]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .X(cubev_phi_din0[12]));
 sky130_fd_sc_hd__clkbuf_4 output396 (.A(net396),
    .X(cubev_phi_din0[13]));
 sky130_fd_sc_hd__clkbuf_4 output397 (.A(net397),
    .X(cubev_phi_din0[14]));
 sky130_fd_sc_hd__clkbuf_4 output398 (.A(net398),
    .X(cubev_phi_din0[15]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .X(cubev_phi_din0[16]));
 sky130_fd_sc_hd__clkbuf_4 output400 (.A(net400),
    .X(cubev_phi_din0[17]));
 sky130_fd_sc_hd__clkbuf_4 output401 (.A(net401),
    .X(cubev_phi_din0[18]));
 sky130_fd_sc_hd__clkbuf_4 output402 (.A(net402),
    .X(cubev_phi_din0[19]));
 sky130_fd_sc_hd__clkbuf_4 output403 (.A(net403),
    .X(cubev_phi_din0[1]));
 sky130_fd_sc_hd__clkbuf_4 output404 (.A(net404),
    .X(cubev_phi_din0[20]));
 sky130_fd_sc_hd__clkbuf_4 output405 (.A(net405),
    .X(cubev_phi_din0[21]));
 sky130_fd_sc_hd__clkbuf_4 output406 (.A(net406),
    .X(cubev_phi_din0[22]));
 sky130_fd_sc_hd__clkbuf_4 output407 (.A(net407),
    .X(cubev_phi_din0[23]));
 sky130_fd_sc_hd__clkbuf_4 output408 (.A(net408),
    .X(cubev_phi_din0[24]));
 sky130_fd_sc_hd__clkbuf_4 output409 (.A(net409),
    .X(cubev_phi_din0[25]));
 sky130_fd_sc_hd__clkbuf_4 output410 (.A(net410),
    .X(cubev_phi_din0[26]));
 sky130_fd_sc_hd__clkbuf_4 output411 (.A(net411),
    .X(cubev_phi_din0[27]));
 sky130_fd_sc_hd__clkbuf_4 output412 (.A(net412),
    .X(cubev_phi_din0[28]));
 sky130_fd_sc_hd__clkbuf_4 output413 (.A(net413),
    .X(cubev_phi_din0[29]));
 sky130_fd_sc_hd__clkbuf_4 output414 (.A(net414),
    .X(cubev_phi_din0[2]));
 sky130_fd_sc_hd__clkbuf_4 output415 (.A(net415),
    .X(cubev_phi_din0[30]));
 sky130_fd_sc_hd__clkbuf_4 output416 (.A(net416),
    .X(cubev_phi_din0[31]));
 sky130_fd_sc_hd__clkbuf_4 output417 (.A(net417),
    .X(cubev_phi_din0[3]));
 sky130_fd_sc_hd__clkbuf_4 output418 (.A(net418),
    .X(cubev_phi_din0[4]));
 sky130_fd_sc_hd__clkbuf_4 output419 (.A(net419),
    .X(cubev_phi_din0[5]));
 sky130_fd_sc_hd__clkbuf_4 output420 (.A(net420),
    .X(cubev_phi_din0[6]));
 sky130_fd_sc_hd__clkbuf_4 output421 (.A(net421),
    .X(cubev_phi_din0[7]));
 sky130_fd_sc_hd__clkbuf_4 output422 (.A(net422),
    .X(cubev_phi_din0[8]));
 sky130_fd_sc_hd__clkbuf_4 output423 (.A(net423),
    .X(cubev_phi_din0[9]));
 sky130_fd_sc_hd__clkbuf_4 output424 (.A(net424),
    .X(cubev_phi_web0));
 sky130_fd_sc_hd__clkbuf_4 output425 (.A(net425),
    .X(cubev_pli_addr0[0]));
 sky130_fd_sc_hd__clkbuf_4 output426 (.A(net426),
    .X(cubev_pli_addr0[1]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .X(cubev_pli_addr0[2]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .X(cubev_pli_addr0[3]));
 sky130_fd_sc_hd__clkbuf_4 output429 (.A(net429),
    .X(cubev_pli_addr0[4]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .X(cubev_pli_addr0[5]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .X(cubev_pli_addr0[6]));
 sky130_fd_sc_hd__clkbuf_4 output432 (.A(net432),
    .X(cubev_pli_addr0[7]));
 sky130_fd_sc_hd__clkbuf_1 output433 (.A(net433),
    .X(cubev_pli_clk0));
 sky130_fd_sc_hd__clkbuf_4 output434 (.A(net434),
    .X(cubev_pli_din0[0]));
 sky130_fd_sc_hd__clkbuf_4 output435 (.A(net435),
    .X(cubev_pli_din0[10]));
 sky130_fd_sc_hd__clkbuf_4 output436 (.A(net436),
    .X(cubev_pli_din0[11]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .X(cubev_pli_din0[12]));
 sky130_fd_sc_hd__clkbuf_4 output438 (.A(net438),
    .X(cubev_pli_din0[13]));
 sky130_fd_sc_hd__clkbuf_4 output439 (.A(net439),
    .X(cubev_pli_din0[14]));
 sky130_fd_sc_hd__clkbuf_4 output440 (.A(net440),
    .X(cubev_pli_din0[15]));
 sky130_fd_sc_hd__clkbuf_4 output441 (.A(net441),
    .X(cubev_pli_din0[16]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .X(cubev_pli_din0[17]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .X(cubev_pli_din0[18]));
 sky130_fd_sc_hd__clkbuf_4 output444 (.A(net444),
    .X(cubev_pli_din0[19]));
 sky130_fd_sc_hd__clkbuf_4 output445 (.A(net445),
    .X(cubev_pli_din0[1]));
 sky130_fd_sc_hd__clkbuf_4 output446 (.A(net446),
    .X(cubev_pli_din0[20]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .X(cubev_pli_din0[21]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .X(cubev_pli_din0[22]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .X(cubev_pli_din0[23]));
 sky130_fd_sc_hd__clkbuf_4 output450 (.A(net450),
    .X(cubev_pli_din0[24]));
 sky130_fd_sc_hd__clkbuf_4 output451 (.A(net451),
    .X(cubev_pli_din0[25]));
 sky130_fd_sc_hd__clkbuf_4 output452 (.A(net452),
    .X(cubev_pli_din0[26]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .X(cubev_pli_din0[27]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .X(cubev_pli_din0[28]));
 sky130_fd_sc_hd__clkbuf_4 output455 (.A(net455),
    .X(cubev_pli_din0[29]));
 sky130_fd_sc_hd__clkbuf_4 output456 (.A(net456),
    .X(cubev_pli_din0[2]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .X(cubev_pli_din0[30]));
 sky130_fd_sc_hd__clkbuf_4 output458 (.A(net458),
    .X(cubev_pli_din0[31]));
 sky130_fd_sc_hd__clkbuf_4 output459 (.A(net459),
    .X(cubev_pli_din0[3]));
 sky130_fd_sc_hd__clkbuf_4 output460 (.A(net460),
    .X(cubev_pli_din0[4]));
 sky130_fd_sc_hd__clkbuf_4 output461 (.A(net461),
    .X(cubev_pli_din0[5]));
 sky130_fd_sc_hd__clkbuf_4 output462 (.A(net462),
    .X(cubev_pli_din0[6]));
 sky130_fd_sc_hd__clkbuf_4 output463 (.A(net463),
    .X(cubev_pli_din0[7]));
 sky130_fd_sc_hd__clkbuf_4 output464 (.A(net464),
    .X(cubev_pli_din0[8]));
 sky130_fd_sc_hd__clkbuf_4 output465 (.A(net465),
    .X(cubev_pli_din0[9]));
 sky130_fd_sc_hd__clkbuf_4 output466 (.A(net466),
    .X(cubev_pli_web0));
 sky130_fd_sc_hd__clkbuf_4 output467 (.A(net467),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output468 (.A(net468),
    .X(la_data_out[100]));
 sky130_fd_sc_hd__clkbuf_4 output469 (.A(net469),
    .X(la_data_out[101]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .X(la_data_out[102]));
 sky130_fd_sc_hd__clkbuf_4 output471 (.A(net471),
    .X(la_data_out[103]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .X(la_data_out[104]));
 sky130_fd_sc_hd__clkbuf_4 output473 (.A(net473),
    .X(la_data_out[105]));
 sky130_fd_sc_hd__clkbuf_4 output474 (.A(net474),
    .X(la_data_out[106]));
 sky130_fd_sc_hd__clkbuf_4 output475 (.A(net475),
    .X(la_data_out[107]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .X(la_data_out[108]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .X(la_data_out[109]));
 sky130_fd_sc_hd__clkbuf_4 output478 (.A(net478),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__clkbuf_4 output479 (.A(net479),
    .X(la_data_out[110]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .X(la_data_out[111]));
 sky130_fd_sc_hd__clkbuf_4 output481 (.A(net481),
    .X(la_data_out[112]));
 sky130_fd_sc_hd__clkbuf_4 output482 (.A(net482),
    .X(la_data_out[113]));
 sky130_fd_sc_hd__clkbuf_4 output483 (.A(net483),
    .X(la_data_out[114]));
 sky130_fd_sc_hd__clkbuf_4 output484 (.A(net484),
    .X(la_data_out[115]));
 sky130_fd_sc_hd__clkbuf_4 output485 (.A(net485),
    .X(la_data_out[116]));
 sky130_fd_sc_hd__clkbuf_4 output486 (.A(net486),
    .X(la_data_out[117]));
 sky130_fd_sc_hd__clkbuf_4 output487 (.A(net487),
    .X(la_data_out[118]));
 sky130_fd_sc_hd__clkbuf_4 output488 (.A(net488),
    .X(la_data_out[119]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__clkbuf_4 output490 (.A(net490),
    .X(la_data_out[120]));
 sky130_fd_sc_hd__clkbuf_4 output491 (.A(net491),
    .X(la_data_out[121]));
 sky130_fd_sc_hd__clkbuf_4 output492 (.A(net492),
    .X(la_data_out[122]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .X(la_data_out[123]));
 sky130_fd_sc_hd__clkbuf_4 output494 (.A(net494),
    .X(la_data_out[124]));
 sky130_fd_sc_hd__clkbuf_4 output495 (.A(net495),
    .X(la_data_out[125]));
 sky130_fd_sc_hd__clkbuf_4 output496 (.A(net496),
    .X(la_data_out[126]));
 sky130_fd_sc_hd__clkbuf_4 output497 (.A(net497),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__clkbuf_4 output498 (.A(net498),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__clkbuf_4 output500 (.A(net500),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__clkbuf_4 output501 (.A(net501),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__clkbuf_4 output502 (.A(net502),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__clkbuf_4 output503 (.A(net503),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__clkbuf_4 output504 (.A(net504),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__clkbuf_4 output505 (.A(net505),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output506 (.A(net506),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__clkbuf_4 output507 (.A(net507),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__clkbuf_4 output508 (.A(net508),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__clkbuf_4 output509 (.A(net509),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__clkbuf_4 output510 (.A(net510),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__clkbuf_4 output511 (.A(net511),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__clkbuf_4 output512 (.A(net512),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__clkbuf_4 output513 (.A(net513),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__clkbuf_4 output514 (.A(net514),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__clkbuf_4 output515 (.A(net515),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__clkbuf_4 output516 (.A(net516),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output517 (.A(net517),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__clkbuf_4 output518 (.A(net518),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__clkbuf_4 output519 (.A(net519),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__clkbuf_4 output520 (.A(net520),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__clkbuf_4 output521 (.A(net521),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__clkbuf_4 output522 (.A(net522),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__clkbuf_4 output523 (.A(net523),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__clkbuf_4 output524 (.A(net524),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__clkbuf_4 output525 (.A(net525),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__clkbuf_4 output526 (.A(net526),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__clkbuf_4 output527 (.A(net527),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__clkbuf_4 output528 (.A(net528),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__clkbuf_4 output529 (.A(net529),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__clkbuf_4 output530 (.A(net530),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__clkbuf_4 output531 (.A(net531),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__clkbuf_4 output532 (.A(net532),
    .X(la_data_out[44]));
 sky130_fd_sc_hd__clkbuf_4 output533 (.A(net533),
    .X(la_data_out[45]));
 sky130_fd_sc_hd__clkbuf_4 output534 (.A(net534),
    .X(la_data_out[46]));
 sky130_fd_sc_hd__clkbuf_4 output535 (.A(net535),
    .X(la_data_out[47]));
 sky130_fd_sc_hd__clkbuf_4 output536 (.A(net536),
    .X(la_data_out[48]));
 sky130_fd_sc_hd__clkbuf_4 output537 (.A(net537),
    .X(la_data_out[49]));
 sky130_fd_sc_hd__clkbuf_4 output538 (.A(net538),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output539 (.A(net539),
    .X(la_data_out[50]));
 sky130_fd_sc_hd__clkbuf_4 output540 (.A(net540),
    .X(la_data_out[51]));
 sky130_fd_sc_hd__clkbuf_4 output541 (.A(net541),
    .X(la_data_out[52]));
 sky130_fd_sc_hd__clkbuf_4 output542 (.A(net542),
    .X(la_data_out[53]));
 sky130_fd_sc_hd__clkbuf_4 output543 (.A(net543),
    .X(la_data_out[54]));
 sky130_fd_sc_hd__clkbuf_4 output544 (.A(net544),
    .X(la_data_out[55]));
 sky130_fd_sc_hd__clkbuf_4 output545 (.A(net545),
    .X(la_data_out[56]));
 sky130_fd_sc_hd__clkbuf_4 output546 (.A(net546),
    .X(la_data_out[57]));
 sky130_fd_sc_hd__clkbuf_4 output547 (.A(net547),
    .X(la_data_out[58]));
 sky130_fd_sc_hd__clkbuf_4 output548 (.A(net548),
    .X(la_data_out[59]));
 sky130_fd_sc_hd__clkbuf_4 output549 (.A(net549),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output550 (.A(net550),
    .X(la_data_out[60]));
 sky130_fd_sc_hd__clkbuf_4 output551 (.A(net551),
    .X(la_data_out[61]));
 sky130_fd_sc_hd__clkbuf_4 output552 (.A(net552),
    .X(la_data_out[62]));
 sky130_fd_sc_hd__clkbuf_4 output553 (.A(net553),
    .X(la_data_out[63]));
 sky130_fd_sc_hd__clkbuf_4 output554 (.A(net554),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__clkbuf_4 output555 (.A(net555),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output556 (.A(net556),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__clkbuf_4 output557 (.A(net557),
    .X(la_data_out[95]));
 sky130_fd_sc_hd__clkbuf_4 output558 (.A(net558),
    .X(la_data_out[96]));
 sky130_fd_sc_hd__clkbuf_4 output559 (.A(net559),
    .X(la_data_out[97]));
 sky130_fd_sc_hd__clkbuf_4 output560 (.A(net560),
    .X(la_data_out[98]));
 sky130_fd_sc_hd__clkbuf_4 output561 (.A(net561),
    .X(la_data_out[99]));
 sky130_fd_sc_hd__clkbuf_4 output562 (.A(net562),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__buf_8 output563 (.A(net630),
    .X(rstn_reg));
 sky130_fd_sc_hd__clkbuf_4 output564 (.A(net564),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__clkbuf_4 output565 (.A(net565),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__clkbuf_4 output566 (.A(net566),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__clkbuf_4 output567 (.A(net567),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__clkbuf_4 output568 (.A(net568),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__clkbuf_4 output569 (.A(net569),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__clkbuf_4 output570 (.A(net570),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__clkbuf_4 output571 (.A(net571),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__clkbuf_4 output572 (.A(net572),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__clkbuf_4 output573 (.A(net573),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__clkbuf_4 output574 (.A(net574),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__clkbuf_4 output575 (.A(net575),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__clkbuf_4 output576 (.A(net576),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__clkbuf_4 output577 (.A(net577),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__clkbuf_4 output578 (.A(net578),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__clkbuf_4 output579 (.A(net579),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__clkbuf_4 output580 (.A(net580),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__clkbuf_4 output581 (.A(net581),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output582 (.A(net582),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output583 (.A(net583),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output584 (.A(net584),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__clkbuf_4 output585 (.A(net585),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__clkbuf_4 output586 (.A(net586),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__clkbuf_4 output587 (.A(net587),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__clkbuf_4 output588 (.A(net588),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__clkbuf_4 output589 (.A(net589),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__clkbuf_4 output590 (.A(net590),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__clkbuf_4 output591 (.A(net591),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__clkbuf_4 output592 (.A(net592),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__clkbuf_4 output593 (.A(net593),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__clkbuf_4 output594 (.A(net594),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__clkbuf_4 output595 (.A(net595),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__clkbuf_8 fanout596 (.A(net602),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_8 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__buf_2 fanout598 (.A(net602),
    .X(net598));
 sky130_fd_sc_hd__buf_6 fanout599 (.A(net601),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_8 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__buf_2 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_6 fanout602 (.A(net563),
    .X(net602));
 sky130_fd_sc_hd__buf_4 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__buf_6 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__buf_6 fanout607 (.A(net632),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_6 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__buf_6 fanout610 (.A(net632),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_4 fanout611 (.A(net632),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_8 fanout612 (.A(net614),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_4 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_8 fanout614 (.A(net623),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__buf_6 fanout616 (.A(net623),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_8 fanout617 (.A(net622),
    .X(net617));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net622),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_8 fanout619 (.A(net622),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_8 fanout620 (.A(net622),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_8 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_6 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(net632),
    .X(net623));
 sky130_fd_sc_hd__buf_6 fanout624 (.A(net626),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_6 fanout626 (.A(net632),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_8 fanout627 (.A(net628),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(net631),
    .X(net628));
 sky130_fd_sc_hd__buf_6 fanout629 (.A(net631),
    .X(net629));
 sky130_fd_sc_hd__buf_8 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__buf_12 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__buf_12 fanout632 (.A(net563),
    .X(net632));
 sky130_fd_sc_hd__conb_1 cawb_633 (.LO(net633));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_opt_5_0_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_wb_clk_i (.A(clknet_1_0_0_wb_clk_i),
    .X(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_wb_clk_i (.A(clknet_1_1_0_wb_clk_i),
    .X(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.A(clknet_1_0_1_wb_clk_i),
    .X(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.A(clknet_1_1_1_wb_clk_i),
    .X(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_opt_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.A(clknet_2_0_0_wb_clk_i),
    .X(clknet_opt_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_1_wb_clk_i (.A(clknet_opt_2_0_wb_clk_i),
    .X(clknet_opt_2_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_2_wb_clk_i (.A(clknet_opt_2_1_wb_clk_i),
    .X(clknet_opt_2_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_3_wb_clk_i (.A(clknet_opt_2_2_wb_clk_i),
    .X(clknet_opt_2_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.A(clknet_2_1_0_wb_clk_i),
    .X(clknet_opt_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_1_wb_clk_i (.A(clknet_opt_3_0_wb_clk_i),
    .X(clknet_opt_3_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_2_wb_clk_i (.A(clknet_opt_3_1_wb_clk_i),
    .X(clknet_opt_3_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_wb_clk_i (.A(clknet_2_2_0_wb_clk_i),
    .X(clknet_opt_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_1_wb_clk_i (.A(clknet_opt_4_0_wb_clk_i),
    .X(clknet_opt_4_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_0_wb_clk_i (.A(clknet_2_3_0_wb_clk_i),
    .X(clknet_opt_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0983_ (.A(_0983_),
    .X(clknet_0__0983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0983_ (.A(clknet_0__0983_),
    .X(clknet_1_0__leaf__0983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0983_ (.A(clknet_0__0983_),
    .X(clknet_1_1__leaf__0983_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1029_ (.A(_1029_),
    .X(clknet_0__1029_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1029_ (.A(clknet_0__1029_),
    .X(clknet_1_0__leaf__1029_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1029_ (.A(clknet_0__1029_),
    .X(clknet_1_1__leaf__1029_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1028_ (.A(_1028_),
    .X(clknet_0__1028_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1028_ (.A(clknet_0__1028_),
    .X(clknet_1_0__leaf__1028_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1028_ (.A(clknet_0__1028_),
    .X(clknet_1_1__leaf__1028_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1027_ (.A(_1027_),
    .X(clknet_0__1027_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1027_ (.A(clknet_0__1027_),
    .X(clknet_1_0__leaf__1027_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1027_ (.A(clknet_0__1027_),
    .X(clknet_1_1__leaf__1027_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1026_ (.A(_1026_),
    .X(clknet_0__1026_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1026_ (.A(clknet_0__1026_),
    .X(clknet_1_0__leaf__1026_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1026_ (.A(clknet_0__1026_),
    .X(clknet_1_1__leaf__1026_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1025_ (.A(_1025_),
    .X(clknet_0__1025_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1025_ (.A(clknet_0__1025_),
    .X(clknet_1_0__leaf__1025_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1025_ (.A(clknet_0__1025_),
    .X(clknet_1_1__leaf__1025_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1024_ (.A(_1024_),
    .X(clknet_0__1024_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1024_ (.A(clknet_0__1024_),
    .X(clknet_1_0__leaf__1024_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1024_ (.A(clknet_0__1024_),
    .X(clknet_1_1__leaf__1024_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0987_ (.A(_0987_),
    .X(clknet_0__0987_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0__0987_ (.A(clknet_0__0987_),
    .X(clknet_1_0_0__0987_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0__0987_ (.A(clknet_0__0987_),
    .X(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1023_ (.A(_1023_),
    .X(clknet_0__1023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1023_ (.A(clknet_0__1023_),
    .X(clknet_1_0__leaf__1023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1023_ (.A(clknet_0__1023_),
    .X(clknet_1_1__leaf__1023_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1022_ (.A(_1022_),
    .X(clknet_0__1022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1022_ (.A(clknet_0__1022_),
    .X(clknet_1_0__leaf__1022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1022_ (.A(clknet_0__1022_),
    .X(clknet_1_1__leaf__1022_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__1021_ (.A(_1021_),
    .X(clknet_0__1021_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__1021_ (.A(clknet_0__1021_),
    .X(clknet_1_0__leaf__1021_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__1021_ (.A(clknet_0__1021_),
    .X(clknet_1_1__leaf__1021_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0994_ (.A(_0994_),
    .X(clknet_0__0994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0994_ (.A(clknet_0__0994_),
    .X(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0994_ (.A(clknet_0__0994_),
    .X(clknet_1_1__leaf__0994_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0993_ (.A(_0993_),
    .X(clknet_0__0993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0993_ (.A(clknet_0__0993_),
    .X(clknet_1_0__leaf__0993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0993_ (.A(clknet_0__0993_),
    .X(clknet_1_1__leaf__0993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0992_ (.A(_0992_),
    .X(clknet_0__0992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0992_ (.A(clknet_0__0992_),
    .X(clknet_1_0__leaf__0992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0992_ (.A(clknet_0__0992_),
    .X(clknet_1_1__leaf__0992_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0991_ (.A(_0991_),
    .X(clknet_0__0991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0991_ (.A(clknet_0__0991_),
    .X(clknet_1_0__leaf__0991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0991_ (.A(clknet_0__0991_),
    .X(clknet_1_1__leaf__0991_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0990_ (.A(_0990_),
    .X(clknet_0__0990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0990_ (.A(clknet_0__0990_),
    .X(clknet_1_0__leaf__0990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0990_ (.A(clknet_0__0990_),
    .X(clknet_1_1__leaf__0990_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0989_ (.A(_0989_),
    .X(clknet_0__0989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0989_ (.A(clknet_0__0989_),
    .X(clknet_1_0__leaf__0989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0989_ (.A(clknet_0__0989_),
    .X(clknet_1_1__leaf__0989_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0988_ (.A(_0988_),
    .X(clknet_0__0988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0988_ (.A(clknet_0__0988_),
    .X(clknet_1_0__leaf__0988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0988_ (.A(clknet_0__0988_),
    .X(clknet_1_1__leaf__0988_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0984_ (.A(_0984_),
    .X(clknet_0__0984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0984_ (.A(clknet_0__0984_),
    .X(clknet_1_0__leaf__0984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0984_ (.A(clknet_0__0984_),
    .X(clknet_1_1__leaf__0984_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0986_ (.A(_0986_),
    .X(clknet_0__0986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0986_ (.A(clknet_0__0986_),
    .X(clknet_1_0__leaf__0986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0986_ (.A(clknet_0__0986_),
    .X(clknet_1_1__leaf__0986_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0985_ (.A(_0985_),
    .X(clknet_0__0985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0985_ (.A(clknet_0__0985_),
    .X(clknet_1_0__leaf__0985_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0985_ (.A(clknet_0__0985_),
    .X(clknet_1_1__leaf__0985_));
 sky130_fd_sc_hd__bufbuf_16 hold1 (.A(\i_ca.ca_rd_fsm_state[1] ),
    .X(net874));
 sky130_fd_sc_hd__bufbuf_16 hold2 (.A(\i_ca.ca_wr_fsm_state[10] ),
    .X(net875));
 sky130_fd_sc_hd__bufbuf_16 hold3 (.A(\i_ca.ca_rd_doutb[32] ),
    .X(net876));
 sky130_fd_sc_hd__bufbuf_16 hold4 (.A(\i_ca.ca_wr_fsm_state[6] ),
    .X(net877));
 sky130_fd_sc_hd__bufbuf_16 hold5 (.A(\i_ca.ca_wr_fsm_state[8] ),
    .X(net878));
 sky130_fd_sc_hd__bufbuf_16 hold6 (.A(\i_ca.ca_wr_fsm_state[17] ),
    .X(net879));
 sky130_fd_sc_hd__bufbuf_16 hold7 (.A(\i_ca.ca_wr_fsm_state[5] ),
    .X(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__D (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A2 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__B (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__C (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__D (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__S (.DIODE(_0012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__D (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A2 (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__S (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A1 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__S (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A1 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__A2 (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__B2 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__B2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__B (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A1_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__B1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A2_N (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__B2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__B (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__B (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A (.DIODE(_0793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__B1 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__S (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__0987__A (.DIODE(_0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__S (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__C (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A2 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__B1 (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__B (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__B (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A2 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__B (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__S (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A2 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__B (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__B2 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__B (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__B (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A0 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__B2 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__B1 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A1 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A1 (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__B2 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__B (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A2 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A2 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A2 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A2 (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A (.DIODE(_1087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__S (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A3 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__B1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__B1 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A2 (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A1 (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__A1 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A1 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__S (.DIODE(_1223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__B1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__B1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__B_N (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A2 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A2 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A2 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A2 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A2 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__B1 (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__A (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__S (.DIODE(_1248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A2 (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__B1 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__B2 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__B1 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__B1 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__B1 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A3 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A2 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A2 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A2 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A2 (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__S (.DIODE(_1279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__B1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__C1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__C1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__B1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__B1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__C1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__B1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__B1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__B1 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__B (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A2 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A2 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__B1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__B2 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__A2 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__B1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__B1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__B1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__C1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A2 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__B1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__S (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__S (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ca_dbus_com));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(ca_dbus_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(ca_dbus_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(ca_dbus_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(ca_dbus_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(ca_dbus_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(ca_dbus_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(ca_dbus_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(ca_dbus_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(ca_dbus_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(ca_dbus_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(ca_dbus_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(ca_dbus_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(ca_dbus_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(ca_dbus_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(ca_dbus_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(ca_dbus_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(ca_dbus_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(ca_dbus_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(ca_dbus_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(ca_dbus_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(ca_dbus_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(ca_dbus_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(ca_dbus_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(ca_dbus_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(ca_dbus_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(ca_dbus_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(ca_dbus_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(ca_dbus_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(ca_dbus_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(ca_dbus_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(ca_dbus_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(ca_dbus_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(ca_dbus_tid[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(ca_dbus_tid[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(ca_dbus_tid[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(ca_dbus_valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(ca_match_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(ca_time_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(cubev_ca_dout0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(cubev_ca_dout0[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(cubev_ca_dout0[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(cubev_ca_dout0[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(cubev_ca_dout0[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(cubev_ca_dout0[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(cubev_ca_dout0[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(cubev_ca_dout0[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(cubev_ca_dout0[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(cubev_ca_dout0[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(cubev_ca_dout0[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(cubev_ca_dout0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(cubev_ca_dout0[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(cubev_ca_dout0[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(cubev_ca_dout0[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(cubev_ca_dout0[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(cubev_ca_dout0[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(cubev_ca_dout0[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(cubev_ca_dout0[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(cubev_ca_dout0[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(cubev_ca_dout0[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(cubev_ca_dout0[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(cubev_ca_dout0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(cubev_ca_dout0[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(cubev_ca_dout0[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(cubev_ca_dout0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(cubev_ca_dout0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(cubev_ca_dout0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(cubev_ca_dout0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(cubev_ca_dout0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(cubev_ca_dout0[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(cubev_ca_dout0[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(cubev_ca_dout1[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(cubev_ca_dout1[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(cubev_ca_dout1[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(cubev_ca_dout1[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(cubev_ca_dout1[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(cubev_ca_dout1[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(cubev_ca_dout1[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(cubev_ca_dout1[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(cubev_ca_dout1[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(cubev_ca_dout1[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(cubev_ca_dout1[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(cubev_ca_dout1[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(cubev_ca_dout1[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(cubev_ca_dout1[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(cubev_ca_dout1[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(cubev_ca_dout1[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(cubev_ca_dout1[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(cubev_ca_dout1[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(cubev_ca_dout1[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(cubev_ca_dout1[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(cubev_ca_dout1[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(cubev_ca_dout1[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(cubev_ca_dout1[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(cubev_ca_dout1[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(cubev_ca_dout1[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(cubev_ca_dout1[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(cubev_ca_dout1[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(cubev_ca_dout1[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(cubev_ca_dout1[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(cubev_ca_dout1[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(cubev_ca_dout1[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(cubev_ca_dout1[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(cubev_phi_dout0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(cubev_phi_dout0[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(cubev_phi_dout0[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(cubev_phi_dout0[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(cubev_phi_dout0[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(cubev_phi_dout0[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(cubev_phi_dout0[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(cubev_phi_dout0[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(cubev_phi_dout0[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(cubev_phi_dout0[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(cubev_phi_dout0[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(cubev_phi_dout0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(cubev_phi_dout0[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(cubev_phi_dout0[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(cubev_phi_dout0[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(cubev_phi_dout0[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(cubev_phi_dout0[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(cubev_phi_dout0[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(cubev_phi_dout0[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(cubev_phi_dout0[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(cubev_phi_dout0[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(cubev_phi_dout0[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(cubev_phi_dout0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(cubev_phi_dout0[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(cubev_phi_dout0[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(cubev_phi_dout0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(cubev_phi_dout0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(cubev_phi_dout0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(cubev_phi_dout0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(cubev_phi_dout0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(cubev_phi_dout0[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(cubev_phi_dout0[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(cubev_pli_dout0[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(cubev_pli_dout0[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(cubev_pli_dout0[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(cubev_pli_dout0[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(cubev_pli_dout0[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(cubev_pli_dout0[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(cubev_pli_dout0[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(cubev_pli_dout0[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(cubev_pli_dout0[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(cubev_pli_dout0[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(cubev_pli_dout0[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(cubev_pli_dout0[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(cubev_pli_dout0[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(cubev_pli_dout0[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(cubev_pli_dout0[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(cubev_pli_dout0[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(cubev_pli_dout0[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(cubev_pli_dout0[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(cubev_pli_dout0[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(cubev_pli_dout0[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(cubev_pli_dout0[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(cubev_pli_dout0[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(cubev_pli_dout0[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(cubev_pli_dout0[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(cubev_pli_dout0[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(cubev_pli_dout0[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(cubev_pli_dout0[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(cubev_pli_dout0[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(cubev_pli_dout0[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(cubev_pli_dout0[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(cubev_pli_dout0[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(cubev_pli_dout0[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A1 (.DIODE(\i_ca.ca_end_of_wr_list ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(\i_ca.ca_end_of_wr_list ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A (.DIODE(\i_ca.ca_end_of_wr_list ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (.DIODE(\i_ca.ca_end_of_wr_list ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A0 (.DIODE(\i_ca.ca_rd_doutb[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A_N (.DIODE(\i_ca.ca_rd_doutb[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A0 (.DIODE(\i_ca.ca_rd_doutb[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__A (.DIODE(\i_ca.ca_rd_doutb[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__B (.DIODE(\i_ca.ca_rd_doutb[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__A0 (.DIODE(\i_ca.ca_rd_doutb[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A1 (.DIODE(\i_ca.ca_rd_doutb[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A1_N (.DIODE(\i_ca.ca_rd_doutb[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__A (.DIODE(\i_ca.ca_rd_doutb[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A0 (.DIODE(\i_ca.ca_rd_doutb[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A (.DIODE(\i_ca.ca_rd_doutb[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__B (.DIODE(\i_ca.ca_rd_doutb[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__C (.DIODE(\i_ca.ca_rd_doutb[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A0 (.DIODE(\i_ca.ca_rd_doutb[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A_N (.DIODE(\i_ca.ca_rd_doutb[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B (.DIODE(\i_ca.ca_rd_doutb[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__B (.DIODE(\i_ca.ca_rd_doutb[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A0 (.DIODE(\i_ca.ca_rd_doutb[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(\i_ca.ca_rd_doutb[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__B_N (.DIODE(\i_ca.ca_rd_doutb[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A (.DIODE(\i_ca.ca_rd_doutb[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A0 (.DIODE(\i_ca.ca_rd_doutb[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__B (.DIODE(\i_ca.ca_rd_doutb[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__A_N (.DIODE(\i_ca.ca_rd_doutb[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__D (.DIODE(\i_ca.ca_rd_doutb[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A0 (.DIODE(\i_ca.ca_rd_doutb[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__B_N (.DIODE(\i_ca.ca_rd_doutb[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__B (.DIODE(\i_ca.ca_rd_doutb[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__C (.DIODE(\i_ca.ca_rd_doutb[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A0 (.DIODE(\i_ca.ca_rd_doutb[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A_N (.DIODE(\i_ca.ca_rd_doutb[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__B (.DIODE(\i_ca.ca_rd_doutb[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__B (.DIODE(\i_ca.ca_rd_doutb[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A0 (.DIODE(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__B1 (.DIODE(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A_N (.DIODE(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__B (.DIODE(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__A (.DIODE(\i_ca.ca_rd_doutb[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A0 (.DIODE(\i_ca.ca_rd_doutb[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A_N (.DIODE(\i_ca.ca_rd_doutb[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__B_N (.DIODE(\i_ca.ca_rd_doutb[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A0 (.DIODE(\i_ca.ca_rd_doutb[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__B (.DIODE(\i_ca.ca_rd_doutb[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__B (.DIODE(\i_ca.ca_rd_doutb[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A0 (.DIODE(\i_ca.ca_rd_doutb[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A2 (.DIODE(\i_ca.ca_rd_doutb[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A (.DIODE(\i_ca.ca_rd_doutb[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A0 (.DIODE(\i_ca.ca_rd_doutb[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A2 (.DIODE(\i_ca.ca_rd_doutb[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__D (.DIODE(\i_ca.ca_rd_doutb[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__A0 (.DIODE(\i_ca.ca_rd_doutb[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A2 (.DIODE(\i_ca.ca_rd_doutb[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__C (.DIODE(\i_ca.ca_rd_doutb[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A0 (.DIODE(\i_ca.ca_rd_doutb[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A2 (.DIODE(\i_ca.ca_rd_doutb[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__B (.DIODE(\i_ca.ca_rd_doutb[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A0 (.DIODE(\i_ca.ca_rd_doutb[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A2 (.DIODE(\i_ca.ca_rd_doutb[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__A (.DIODE(\i_ca.ca_rd_doutb[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A0 (.DIODE(\i_ca.ca_rd_doutb[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A2 (.DIODE(\i_ca.ca_rd_doutb[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__D (.DIODE(\i_ca.ca_rd_doutb[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A0 (.DIODE(\i_ca.ca_rd_doutb[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__A (.DIODE(\i_ca.ca_rd_doutb[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A0 (.DIODE(\i_ca.ca_rd_doutb[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A2 (.DIODE(\i_ca.ca_rd_doutb[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__C (.DIODE(\i_ca.ca_rd_doutb[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A0 (.DIODE(\i_ca.ca_rd_doutb[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A (.DIODE(\i_ca.ca_rd_doutb[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A0 (.DIODE(\i_ca.ca_rd_doutb[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A (.DIODE(\i_ca.ca_rd_doutb[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A0 (.DIODE(\i_ca.ca_rd_doutb[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(\i_ca.ca_rd_doutb[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__A0 (.DIODE(\i_ca.ca_rd_doutb[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A (.DIODE(\i_ca.ca_rd_doutb[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__A0 (.DIODE(\i_ca.ca_rd_doutb[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A (.DIODE(\i_ca.ca_rd_doutb[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A0 (.DIODE(\i_ca.ca_rd_doutb[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A (.DIODE(\i_ca.ca_rd_doutb[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__A0 (.DIODE(\i_ca.ca_rd_doutb[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__A (.DIODE(\i_ca.ca_rd_doutb[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B (.DIODE(\i_ca.ca_rd_doutb[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__B (.DIODE(\i_ca.ca_rd_doutb_32 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A1 (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A_N (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__B (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__A1 (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A_N (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__B (.DIODE(\i_ca.ca_ready ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A1 (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__A (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__B2 (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__B1 (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__A (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__B (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1711__A (.DIODE(\i_ca.ca_update_rd_add ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__D (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A1 (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A1 (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A1 (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__A2 (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A (.DIODE(\i_ca.ca_wr_add[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__D (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A2 (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__B2 (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__B (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__B (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A2 (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__B (.DIODE(\i_ca.ca_wr_add[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__D (.DIODE(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A1 (.DIODE(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__B1 (.DIODE(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__A2 (.DIODE(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__C (.DIODE(\i_ca.ca_wr_add[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__D (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A1 (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A1 (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A2 (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__A (.DIODE(\i_ca.ca_wr_add[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__D (.DIODE(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__B1 (.DIODE(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A2 (.DIODE(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__B (.DIODE(\i_ca.ca_wr_add[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__D (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__B2 (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A2 (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__A (.DIODE(\i_ca.ca_wr_add[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__D (.DIODE(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__B1 (.DIODE(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__B (.DIODE(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A2 (.DIODE(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__B (.DIODE(\i_ca.ca_wr_add[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__D (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__A1 (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A1 (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A2 (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__A (.DIODE(\i_ca.ca_wr_add[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__B2 (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A1 (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A1 (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__B2 (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__A (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__B1 (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__A (.DIODE(\i_ca.ca_wr_add_fill[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A1 (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A1 (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A1 (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__B2 (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__C (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A1 (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__B (.DIODE(\i_ca.ca_wr_add_fill[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__B2 (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A1 (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A1 (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B2 (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A1 (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__B (.DIODE(\i_ca.ca_wr_add_fill[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A1 (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__B2 (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A1 (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A1 (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__B (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__C_N (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__A (.DIODE(\i_ca.ca_wr_add_fill[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A1 (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__B2 (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__A1 (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__B2 (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A1 (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__D_N (.DIODE(\i_ca.ca_wr_add_fill[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B2 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A1 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A1 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__B2 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A2 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A1 (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__B (.DIODE(\i_ca.ca_wr_add_fill[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B2 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__B2 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A1 (.DIODE(\i_ca.ca_wr_add_fill[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__C (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__B2 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__B1 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__C (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__B2 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A0 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__B1 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A1 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__A1 (.DIODE(\i_ca.ca_wr_add_start[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A2 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A1 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__S (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A1 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__B1 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A1 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__A1 (.DIODE(\i_ca.ca_wr_add_start[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__B1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__B (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__B1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__B1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A1 (.DIODE(\i_ca.ca_wr_add_start[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__B (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__A1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A1 (.DIODE(\i_ca.ca_wr_add_start[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A1 (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A1 (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__B1 (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__B1 (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(\i_ca.ca_wr_com_const ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__D (.DIODE(\i_ca.ca_wr_dina[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A2 (.DIODE(\i_ca.ca_wr_dina[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A1 (.DIODE(\i_ca.ca_wr_dina[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__D (.DIODE(\i_ca.ca_wr_dina[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A0 (.DIODE(\i_ca.ca_wr_dina[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A1 (.DIODE(\i_ca.ca_wr_dina[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__D (.DIODE(\i_ca.ca_wr_dina[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A0 (.DIODE(\i_ca.ca_wr_dina[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A1 (.DIODE(\i_ca.ca_wr_dina[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__D (.DIODE(\i_ca.ca_wr_dina[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A0 (.DIODE(\i_ca.ca_wr_dina[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A1 (.DIODE(\i_ca.ca_wr_dina[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__D (.DIODE(\i_ca.ca_wr_dina[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A0 (.DIODE(\i_ca.ca_wr_dina[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A1 (.DIODE(\i_ca.ca_wr_dina[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__D (.DIODE(\i_ca.ca_wr_dina[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A0 (.DIODE(\i_ca.ca_wr_dina[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A1 (.DIODE(\i_ca.ca_wr_dina[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__D (.DIODE(\i_ca.ca_wr_dina[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A0 (.DIODE(\i_ca.ca_wr_dina[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A1 (.DIODE(\i_ca.ca_wr_dina[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__D (.DIODE(\i_ca.ca_wr_dina[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A0 (.DIODE(\i_ca.ca_wr_dina[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A1 (.DIODE(\i_ca.ca_wr_dina[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__D (.DIODE(\i_ca.ca_wr_dina[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A0 (.DIODE(\i_ca.ca_wr_dina[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(\i_ca.ca_wr_douta[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A2 (.DIODE(\i_ca.ca_wr_douta[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__A2 (.DIODE(\i_ca.ca_wr_douta[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__B2 (.DIODE(\i_ca.ca_wr_douta[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A2 (.DIODE(\i_ca.ca_wr_douta[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__A2 (.DIODE(\i_ca.ca_wr_douta[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__B2 (.DIODE(\i_ca.ca_wr_douta[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (.DIODE(\i_ca.ca_wr_douta[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A1 (.DIODE(\i_ca.ca_wr_douta[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A (.DIODE(\i_ca.ca_wr_douta[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__B1 (.DIODE(\i_ca.ca_wr_douta[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A (.DIODE(\i_ca.ca_wr_douta[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A (.DIODE(\i_ca.ca_wr_douta[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A1 (.DIODE(\i_ca.ca_wr_douta[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A (.DIODE(\i_ca.ca_wr_douta[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A1 (.DIODE(\i_ca.ca_wr_douta[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A (.DIODE(\i_ca.ca_wr_douta[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A (.DIODE(\i_ca.ca_wr_douta[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A (.DIODE(\i_ca.ca_wr_douta[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1822__B2 (.DIODE(\i_ca.ca_wr_douta[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__B (.DIODE(\i_ca.ca_wr_douta[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__B2 (.DIODE(\i_ca.ca_wr_douta[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(\i_ca.ca_wr_douta[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__B2 (.DIODE(\i_ca.ca_wr_douta[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__A (.DIODE(\i_ca.ca_wr_douta[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B2 (.DIODE(\i_ca.ca_wr_douta[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A (.DIODE(\i_ca.ca_wr_douta[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__B (.DIODE(\i_ca.ca_wr_douta[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__A3 (.DIODE(\i_ca.ca_wr_douta[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A2 (.DIODE(\i_ca.ca_wr_douta[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__B (.DIODE(\i_ca.ca_wr_douta[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A1 (.DIODE(\i_ca.ca_wr_douta[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A2 (.DIODE(\i_ca.ca_wr_douta[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__A (.DIODE(\i_ca.ca_wr_douta[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A1 (.DIODE(\i_ca.ca_wr_douta[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A2 (.DIODE(\i_ca.ca_wr_douta[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__D (.DIODE(\i_ca.ca_wr_douta[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A (.DIODE(\i_ca.ca_wr_douta[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A2 (.DIODE(\i_ca.ca_wr_douta[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A (.DIODE(\i_ca.ca_wr_douta[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A1 (.DIODE(\i_ca.ca_wr_douta[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A2 (.DIODE(\i_ca.ca_wr_douta[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__C (.DIODE(\i_ca.ca_wr_douta[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__A2 (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A2 (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A1 (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__B (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__A_N (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A2 (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A_N (.DIODE(\i_ca.ca_wr_douta[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A (.DIODE(\i_ca.ca_wr_douta[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__A (.DIODE(\i_ca.ca_wr_douta[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A (.DIODE(\i_ca.ca_wr_douta[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__B (.DIODE(\i_ca.ca_wr_douta[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A2 (.DIODE(\i_ca.ca_wr_douta[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A (.DIODE(\i_ca.ca_wr_douta[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A2 (.DIODE(\i_ca.ca_wr_douta[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__B (.DIODE(\i_ca.ca_wr_douta[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__D (.DIODE(\i_ca.ca_wr_fsm_state[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__C (.DIODE(\i_ca.ca_wr_fsm_state[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A1_N (.DIODE(\i_ca.ca_wr_fsm_state[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__B2 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(\i_ca.hs_write_dbus_wr_data_const[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A2 (.DIODE(\i_ca.hs_write_tid_wr0_const[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__A1 (.DIODE(\i_ca.hs_write_tid_wr0_const[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A1 (.DIODE(\i_ca.hs_write_tid_wr0_const[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A1 (.DIODE(\i_ca.hs_write_tid_wr0_const[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(\i_ca.hs_write_tid_wr0_const[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A1 (.DIODE(\i_ca.hs_write_tid_wr0_const[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(la_data_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(la_data_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(la_data_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(la_data_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(la_data_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(la_data_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(la_data_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(la_data_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(la_data_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(la_data_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(la_data_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(la_data_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(la_data_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(la_data_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(la_data_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(la_data_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(la_data_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(la_data_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(la_data_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(la_data_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(la_data_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(la_data_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(la_data_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(la_data_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(la_data_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(la_data_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(la_data_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(la_data_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(la_data_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(la_data_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(la_data_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input199_A (.DIODE(la_data_in[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input200_A (.DIODE(la_data_in[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input201_A (.DIODE(la_data_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input202_A (.DIODE(la_data_in[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input203_A (.DIODE(la_data_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input204_A (.DIODE(la_data_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input205_A (.DIODE(la_data_in[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input206_A (.DIODE(la_data_in[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input207_A (.DIODE(la_data_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input208_A (.DIODE(la_data_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input209_A (.DIODE(la_data_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input210_A (.DIODE(la_data_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input211_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input212_A (.DIODE(wbs_adr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input213_A (.DIODE(wbs_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input214_A (.DIODE(wbs_adr_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input215_A (.DIODE(wbs_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input216_A (.DIODE(wbs_adr_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input217_A (.DIODE(wbs_adr_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input218_A (.DIODE(wbs_adr_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input219_A (.DIODE(wbs_adr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input220_A (.DIODE(wbs_adr_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input221_A (.DIODE(wbs_adr_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input222_A (.DIODE(wbs_adr_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input223_A (.DIODE(wbs_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input224_A (.DIODE(wbs_adr_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input225_A (.DIODE(wbs_adr_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input226_A (.DIODE(wbs_adr_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input227_A (.DIODE(wbs_adr_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input228_A (.DIODE(wbs_adr_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input229_A (.DIODE(wbs_adr_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input230_A (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input231_A (.DIODE(wbs_adr_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input232_A (.DIODE(wbs_adr_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input233_A (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input234_A (.DIODE(wbs_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input235_A (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input236_A (.DIODE(wbs_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input237_A (.DIODE(wbs_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input238_A (.DIODE(wbs_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input239_A (.DIODE(wbs_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input240_A (.DIODE(wbs_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input241_A (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input242_A (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input243_A (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input244_A (.DIODE(wbs_dat_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input245_A (.DIODE(wbs_dat_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input246_A (.DIODE(wbs_dat_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input247_A (.DIODE(wbs_dat_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input248_A (.DIODE(wbs_dat_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input249_A (.DIODE(wbs_dat_i[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input250_A (.DIODE(wbs_dat_i[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input251_A (.DIODE(wbs_dat_i[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input252_A (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input253_A (.DIODE(wbs_dat_i[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input254_A (.DIODE(wbs_dat_i[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input255_A (.DIODE(wbs_dat_i[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input256_A (.DIODE(wbs_dat_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input257_A (.DIODE(wbs_dat_i[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input258_A (.DIODE(wbs_dat_i[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input259_A (.DIODE(wbs_dat_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input260_A (.DIODE(wbs_dat_i[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input261_A (.DIODE(wbs_dat_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input262_A (.DIODE(wbs_dat_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input263_A (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input264_A (.DIODE(wbs_dat_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input265_A (.DIODE(wbs_dat_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input266_A (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input267_A (.DIODE(wbs_dat_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input268_A (.DIODE(wbs_dat_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input269_A (.DIODE(wbs_dat_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input270_A (.DIODE(wbs_dat_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input271_A (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input272_A (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input273_A (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input274_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A0 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__D (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__D (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__D (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__D (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__D (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__D (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__D (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__D (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__D (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__D (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__D (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__D (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__D (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__D (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__D (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__D (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__D (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__D (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__D (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__D (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__D (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__D (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__D (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__D (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__D (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__D (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__D (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__D (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__D (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__D (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__D (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__D (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__B (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__D (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__D (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__D (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__D (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__D (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__D (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__D (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__D (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__D (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__D (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__D (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__D (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__D (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__D (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__D (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__D (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__D (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__D (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__D (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__D (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__A1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__D (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__D (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output277_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__D (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_output278_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__D (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_output279_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__D (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_output280_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__D (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__D (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__D (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_output283_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__D (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__D (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_output285_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__D (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_output286_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__D (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_output287_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__D (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__D (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__D (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__D (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__D (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__D (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__D (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__D (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__D (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__D (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__D (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__D (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__D (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__D (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__D (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__D (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__D (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__D (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__D (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output382_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_output383_A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A0 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_output384_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__A0 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_output385_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A0 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_output386_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_output387_A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__A0 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_output388_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A0 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_output389_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__A0 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_output390_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_output392_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__A0 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_output393_A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__A0 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA_output394_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A0 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_output395_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A0 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_output396_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_output397_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A0 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_output399_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A0 (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_output400_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_output401_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A0 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A0 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_output403_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A0 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_output404_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A0 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A0 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A0 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A0 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_output410_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A0 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_output411_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A0 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A0 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_output413_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A0 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__A0 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__A0 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_output418_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__A0 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__1564__A0 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__A0 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__A0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A0 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A0 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output451_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_output455_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output458_A (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_output482_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_output483_A (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_output484_A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_output485_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_output486_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_output487_A (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_output488_A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_output491_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_output492_A (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_output493_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_output494_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_output495_A (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_output496_A (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_output557_A (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_output573_A (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA_output574_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_output580_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_output582_A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_output587_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_output588_A (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout598_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__B1 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__RESET_B (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__RESET_B (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__RESET_B (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__RESET_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__RESET_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__RESET_B (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__RESET_B (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__RESET_B (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__RESET_B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__RESET_B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__RESET_B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__RESET_B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__RESET_B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__SET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__RESET_B (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__RESET_B (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__RESET_B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__RESET_B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__RESET_B (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__RESET_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__RESET_B (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__RESET_B (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__RESET_B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__RESET_B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout630_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__RESET_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__RESET_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__RESET_B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout631_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_wb_clk_i_A (.DIODE(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_wb_clk_i_A (.DIODE(clknet_1_0_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_wb_clk_i_A (.DIODE(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_wb_clk_i_A (.DIODE(clknet_1_1_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_3_0_wb_clk_i_A (.DIODE(clknet_2_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_4_0_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_2_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_5_0_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_3_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__A (.DIODE(clknet_opt_1_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A (.DIODE(clknet_opt_2_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A (.DIODE(clknet_opt_3_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0__0987__A (.DIODE(clknet_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0__0987__A (.DIODE(clknet_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A (.DIODE(clknet_1_0_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A (.DIODE(clknet_1_0_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__A (.DIODE(clknet_1_0_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A (.DIODE(clknet_1_0_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(clknet_1_1_0__0987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__153_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__154_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__155_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__156_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__157_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__158_A (.DIODE(clknet_1_0__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__149_A (.DIODE(clknet_1_1__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__150_A (.DIODE(clknet_1_1__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__151_A (.DIODE(clknet_1_1__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__152_A (.DIODE(clknet_1_1__leaf__0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__A (.DIODE(clknet_1_1__leaf__0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A (.DIODE(clknet_1_1__leaf__0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__1_A (.DIODE(clknet_1_1__leaf__0984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__8_A (.DIODE(clknet_1_1__leaf__0984_));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1055 ();
 assign ca_command[31] = net633;
 assign cubev_ca_csb0 = net634;
 assign cubev_ca_csb1 = net635;
 assign cubev_ca_wmask0[0] = net674;
 assign cubev_ca_wmask0[1] = net675;
 assign cubev_ca_wmask0[2] = net676;
 assign cubev_ca_wmask0[3] = net677;
 assign cubev_phi_csb0 = net636;
 assign cubev_phi_wmask0[0] = net678;
 assign cubev_phi_wmask0[1] = net679;
 assign cubev_phi_wmask0[2] = net680;
 assign cubev_phi_wmask0[3] = net681;
 assign cubev_pli_csb0 = net637;
 assign cubev_pli_wmask0[0] = net682;
 assign cubev_pli_wmask0[1] = net683;
 assign cubev_pli_wmask0[2] = net684;
 assign cubev_pli_wmask0[3] = net685;
 assign irq[0] = net638;
 assign irq[1] = net639;
 assign irq[2] = net640;
 assign la_data_out[127] = net672;
 assign la_data_out[64] = net641;
 assign la_data_out[65] = net642;
 assign la_data_out[66] = net643;
 assign la_data_out[67] = net644;
 assign la_data_out[68] = net645;
 assign la_data_out[69] = net646;
 assign la_data_out[70] = net647;
 assign la_data_out[71] = net648;
 assign la_data_out[72] = net649;
 assign la_data_out[73] = net650;
 assign la_data_out[74] = net651;
 assign la_data_out[75] = net652;
 assign la_data_out[76] = net653;
 assign la_data_out[77] = net654;
 assign la_data_out[78] = net655;
 assign la_data_out[79] = net656;
 assign la_data_out[80] = net657;
 assign la_data_out[81] = net658;
 assign la_data_out[82] = net659;
 assign la_data_out[83] = net660;
 assign la_data_out[84] = net661;
 assign la_data_out[85] = net662;
 assign la_data_out[86] = net663;
 assign la_data_out[87] = net664;
 assign la_data_out[88] = net665;
 assign la_data_out[89] = net666;
 assign la_data_out[90] = net667;
 assign la_data_out[91] = net668;
 assign la_data_out[92] = net669;
 assign la_data_out[93] = net670;
 assign la_data_out[94] = net671;
 assign wbs_ack_o = net673;
endmodule

