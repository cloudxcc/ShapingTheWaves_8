VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cawb
  CLASS BLOCK ;
  FOREIGN cawb ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 400.000 ;
  PIN ca_command[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 396.000 404.710 400.000 ;
    END
  END ca_command[0]
  PIN ca_command[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 396.000 432.310 400.000 ;
    END
  END ca_command[10]
  PIN ca_command[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 396.000 435.070 400.000 ;
    END
  END ca_command[11]
  PIN ca_command[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 396.000 437.830 400.000 ;
    END
  END ca_command[12]
  PIN ca_command[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 396.000 440.590 400.000 ;
    END
  END ca_command[13]
  PIN ca_command[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 396.000 443.350 400.000 ;
    END
  END ca_command[14]
  PIN ca_command[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 396.000 446.110 400.000 ;
    END
  END ca_command[15]
  PIN ca_command[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 396.000 448.870 400.000 ;
    END
  END ca_command[16]
  PIN ca_command[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 396.000 451.630 400.000 ;
    END
  END ca_command[17]
  PIN ca_command[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 396.000 454.390 400.000 ;
    END
  END ca_command[18]
  PIN ca_command[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 396.000 457.150 400.000 ;
    END
  END ca_command[19]
  PIN ca_command[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 396.000 407.470 400.000 ;
    END
  END ca_command[1]
  PIN ca_command[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 396.000 459.910 400.000 ;
    END
  END ca_command[20]
  PIN ca_command[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 396.000 462.670 400.000 ;
    END
  END ca_command[21]
  PIN ca_command[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 396.000 465.430 400.000 ;
    END
  END ca_command[22]
  PIN ca_command[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 396.000 468.190 400.000 ;
    END
  END ca_command[23]
  PIN ca_command[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 396.000 470.950 400.000 ;
    END
  END ca_command[24]
  PIN ca_command[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 396.000 473.710 400.000 ;
    END
  END ca_command[25]
  PIN ca_command[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 396.000 476.470 400.000 ;
    END
  END ca_command[26]
  PIN ca_command[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 396.000 479.230 400.000 ;
    END
  END ca_command[27]
  PIN ca_command[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 396.000 481.990 400.000 ;
    END
  END ca_command[28]
  PIN ca_command[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 396.000 484.750 400.000 ;
    END
  END ca_command[29]
  PIN ca_command[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 396.000 410.230 400.000 ;
    END
  END ca_command[2]
  PIN ca_command[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 396.000 487.510 400.000 ;
    END
  END ca_command[30]
  PIN ca_command[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 396.000 490.270 400.000 ;
    END
  END ca_command[31]
  PIN ca_command[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 396.000 412.990 400.000 ;
    END
  END ca_command[3]
  PIN ca_command[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 396.000 415.750 400.000 ;
    END
  END ca_command[4]
  PIN ca_command[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 396.000 418.510 400.000 ;
    END
  END ca_command[5]
  PIN ca_command[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 396.000 421.270 400.000 ;
    END
  END ca_command[6]
  PIN ca_command[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 396.000 424.030 400.000 ;
    END
  END ca_command[7]
  PIN ca_command[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 396.000 426.790 400.000 ;
    END
  END ca_command[8]
  PIN ca_command[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 396.000 429.550 400.000 ;
    END
  END ca_command[9]
  PIN ca_dbus_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 396.000 228.070 400.000 ;
    END
  END ca_dbus_ack
  PIN ca_dbus_com
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 396.000 230.830 400.000 ;
    END
  END ca_dbus_com
  PIN ca_dbus_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 396.000 241.870 400.000 ;
    END
  END ca_dbus_data[0]
  PIN ca_dbus_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 396.000 269.470 400.000 ;
    END
  END ca_dbus_data[10]
  PIN ca_dbus_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 396.000 272.230 400.000 ;
    END
  END ca_dbus_data[11]
  PIN ca_dbus_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 396.000 274.990 400.000 ;
    END
  END ca_dbus_data[12]
  PIN ca_dbus_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 396.000 277.750 400.000 ;
    END
  END ca_dbus_data[13]
  PIN ca_dbus_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 396.000 280.510 400.000 ;
    END
  END ca_dbus_data[14]
  PIN ca_dbus_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 396.000 283.270 400.000 ;
    END
  END ca_dbus_data[15]
  PIN ca_dbus_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 396.000 286.030 400.000 ;
    END
  END ca_dbus_data[16]
  PIN ca_dbus_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 396.000 288.790 400.000 ;
    END
  END ca_dbus_data[17]
  PIN ca_dbus_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 396.000 291.550 400.000 ;
    END
  END ca_dbus_data[18]
  PIN ca_dbus_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 396.000 294.310 400.000 ;
    END
  END ca_dbus_data[19]
  PIN ca_dbus_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 396.000 244.630 400.000 ;
    END
  END ca_dbus_data[1]
  PIN ca_dbus_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 396.000 297.070 400.000 ;
    END
  END ca_dbus_data[20]
  PIN ca_dbus_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 396.000 299.830 400.000 ;
    END
  END ca_dbus_data[21]
  PIN ca_dbus_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 396.000 302.590 400.000 ;
    END
  END ca_dbus_data[22]
  PIN ca_dbus_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 396.000 305.350 400.000 ;
    END
  END ca_dbus_data[23]
  PIN ca_dbus_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 396.000 308.110 400.000 ;
    END
  END ca_dbus_data[24]
  PIN ca_dbus_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 396.000 310.870 400.000 ;
    END
  END ca_dbus_data[25]
  PIN ca_dbus_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 396.000 313.630 400.000 ;
    END
  END ca_dbus_data[26]
  PIN ca_dbus_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 396.000 316.390 400.000 ;
    END
  END ca_dbus_data[27]
  PIN ca_dbus_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 396.000 319.150 400.000 ;
    END
  END ca_dbus_data[28]
  PIN ca_dbus_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 396.000 321.910 400.000 ;
    END
  END ca_dbus_data[29]
  PIN ca_dbus_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 396.000 247.390 400.000 ;
    END
  END ca_dbus_data[2]
  PIN ca_dbus_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 396.000 324.670 400.000 ;
    END
  END ca_dbus_data[30]
  PIN ca_dbus_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 396.000 327.430 400.000 ;
    END
  END ca_dbus_data[31]
  PIN ca_dbus_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 396.000 250.150 400.000 ;
    END
  END ca_dbus_data[3]
  PIN ca_dbus_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 396.000 252.910 400.000 ;
    END
  END ca_dbus_data[4]
  PIN ca_dbus_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 396.000 255.670 400.000 ;
    END
  END ca_dbus_data[5]
  PIN ca_dbus_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 396.000 258.430 400.000 ;
    END
  END ca_dbus_data[6]
  PIN ca_dbus_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 396.000 261.190 400.000 ;
    END
  END ca_dbus_data[7]
  PIN ca_dbus_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 396.000 263.950 400.000 ;
    END
  END ca_dbus_data[8]
  PIN ca_dbus_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 396.000 266.710 400.000 ;
    END
  END ca_dbus_data[9]
  PIN ca_dbus_tid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 396.000 233.590 400.000 ;
    END
  END ca_dbus_tid[0]
  PIN ca_dbus_tid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 396.000 236.350 400.000 ;
    END
  END ca_dbus_tid[1]
  PIN ca_dbus_tid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 396.000 239.110 400.000 ;
    END
  END ca_dbus_tid[2]
  PIN ca_dbus_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 396.000 225.310 400.000 ;
    END
  END ca_dbus_valid
  PIN ca_match_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 396.000 401.950 400.000 ;
    END
  END ca_match_ack
  PIN ca_match_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 396.000 399.190 400.000 ;
    END
  END ca_match_valid
  PIN ca_time_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 396.000 332.950 400.000 ;
    END
  END ca_time_ack
  PIN ca_time_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 396.000 335.710 400.000 ;
    END
  END ca_time_data[0]
  PIN ca_time_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 396.000 363.310 400.000 ;
    END
  END ca_time_data[10]
  PIN ca_time_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 396.000 366.070 400.000 ;
    END
  END ca_time_data[11]
  PIN ca_time_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 396.000 368.830 400.000 ;
    END
  END ca_time_data[12]
  PIN ca_time_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 396.000 371.590 400.000 ;
    END
  END ca_time_data[13]
  PIN ca_time_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 396.000 374.350 400.000 ;
    END
  END ca_time_data[14]
  PIN ca_time_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 396.000 377.110 400.000 ;
    END
  END ca_time_data[15]
  PIN ca_time_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 396.000 379.870 400.000 ;
    END
  END ca_time_data[16]
  PIN ca_time_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 396.000 382.630 400.000 ;
    END
  END ca_time_data[17]
  PIN ca_time_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 396.000 385.390 400.000 ;
    END
  END ca_time_data[18]
  PIN ca_time_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 396.000 388.150 400.000 ;
    END
  END ca_time_data[19]
  PIN ca_time_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 396.000 338.470 400.000 ;
    END
  END ca_time_data[1]
  PIN ca_time_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 396.000 390.910 400.000 ;
    END
  END ca_time_data[20]
  PIN ca_time_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 396.000 393.670 400.000 ;
    END
  END ca_time_data[21]
  PIN ca_time_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 396.000 396.430 400.000 ;
    END
  END ca_time_data[22]
  PIN ca_time_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 396.000 341.230 400.000 ;
    END
  END ca_time_data[2]
  PIN ca_time_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 396.000 343.990 400.000 ;
    END
  END ca_time_data[3]
  PIN ca_time_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 396.000 346.750 400.000 ;
    END
  END ca_time_data[4]
  PIN ca_time_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 396.000 349.510 400.000 ;
    END
  END ca_time_data[5]
  PIN ca_time_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END ca_time_data[6]
  PIN ca_time_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 396.000 355.030 400.000 ;
    END
  END ca_time_data[7]
  PIN ca_time_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 396.000 357.790 400.000 ;
    END
  END ca_time_data[8]
  PIN ca_time_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 396.000 360.550 400.000 ;
    END
  END ca_time_data[9]
  PIN ca_time_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 396.000 330.190 400.000 ;
    END
  END ca_time_valid
  PIN cubev_ca_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 55.120 500.000 55.720 ;
    END
  END cubev_ca_addr0[0]
  PIN cubev_ca_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END cubev_ca_addr0[1]
  PIN cubev_ca_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 60.560 500.000 61.160 ;
    END
  END cubev_ca_addr0[2]
  PIN cubev_ca_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 63.280 500.000 63.880 ;
    END
  END cubev_ca_addr0[3]
  PIN cubev_ca_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 66.000 500.000 66.600 ;
    END
  END cubev_ca_addr0[4]
  PIN cubev_ca_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.720 500.000 69.320 ;
    END
  END cubev_ca_addr0[5]
  PIN cubev_ca_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 71.440 500.000 72.040 ;
    END
  END cubev_ca_addr0[6]
  PIN cubev_ca_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 74.160 500.000 74.760 ;
    END
  END cubev_ca_addr0[7]
  PIN cubev_ca_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 256.400 500.000 257.000 ;
    END
  END cubev_ca_addr1[0]
  PIN cubev_ca_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 259.120 500.000 259.720 ;
    END
  END cubev_ca_addr1[1]
  PIN cubev_ca_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 261.840 500.000 262.440 ;
    END
  END cubev_ca_addr1[2]
  PIN cubev_ca_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 264.560 500.000 265.160 ;
    END
  END cubev_ca_addr1[3]
  PIN cubev_ca_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 267.280 500.000 267.880 ;
    END
  END cubev_ca_addr1[4]
  PIN cubev_ca_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 270.000 500.000 270.600 ;
    END
  END cubev_ca_addr1[5]
  PIN cubev_ca_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 272.720 500.000 273.320 ;
    END
  END cubev_ca_addr1[6]
  PIN cubev_ca_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END cubev_ca_addr1[7]
  PIN cubev_ca_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.080 500.000 36.680 ;
    END
  END cubev_ca_clk0
  PIN cubev_ca_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 250.960 500.000 251.560 ;
    END
  END cubev_ca_clk1
  PIN cubev_ca_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 38.800 500.000 39.400 ;
    END
  END cubev_ca_csb0
  PIN cubev_ca_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 253.680 500.000 254.280 ;
    END
  END cubev_ca_csb1
  PIN cubev_ca_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.880 500.000 77.480 ;
    END
  END cubev_ca_din0[0]
  PIN cubev_ca_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 104.080 500.000 104.680 ;
    END
  END cubev_ca_din0[10]
  PIN cubev_ca_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 106.800 500.000 107.400 ;
    END
  END cubev_ca_din0[11]
  PIN cubev_ca_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 109.520 500.000 110.120 ;
    END
  END cubev_ca_din0[12]
  PIN cubev_ca_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END cubev_ca_din0[13]
  PIN cubev_ca_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 114.960 500.000 115.560 ;
    END
  END cubev_ca_din0[14]
  PIN cubev_ca_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 117.680 500.000 118.280 ;
    END
  END cubev_ca_din0[15]
  PIN cubev_ca_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 120.400 500.000 121.000 ;
    END
  END cubev_ca_din0[16]
  PIN cubev_ca_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 123.120 500.000 123.720 ;
    END
  END cubev_ca_din0[17]
  PIN cubev_ca_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 125.840 500.000 126.440 ;
    END
  END cubev_ca_din0[18]
  PIN cubev_ca_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 128.560 500.000 129.160 ;
    END
  END cubev_ca_din0[19]
  PIN cubev_ca_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 79.600 500.000 80.200 ;
    END
  END cubev_ca_din0[1]
  PIN cubev_ca_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 131.280 500.000 131.880 ;
    END
  END cubev_ca_din0[20]
  PIN cubev_ca_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 134.000 500.000 134.600 ;
    END
  END cubev_ca_din0[21]
  PIN cubev_ca_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 136.720 500.000 137.320 ;
    END
  END cubev_ca_din0[22]
  PIN cubev_ca_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 139.440 500.000 140.040 ;
    END
  END cubev_ca_din0[23]
  PIN cubev_ca_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.160 500.000 142.760 ;
    END
  END cubev_ca_din0[24]
  PIN cubev_ca_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 144.880 500.000 145.480 ;
    END
  END cubev_ca_din0[25]
  PIN cubev_ca_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 147.600 500.000 148.200 ;
    END
  END cubev_ca_din0[26]
  PIN cubev_ca_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 150.320 500.000 150.920 ;
    END
  END cubev_ca_din0[27]
  PIN cubev_ca_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 153.040 500.000 153.640 ;
    END
  END cubev_ca_din0[28]
  PIN cubev_ca_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.760 500.000 156.360 ;
    END
  END cubev_ca_din0[29]
  PIN cubev_ca_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 82.320 500.000 82.920 ;
    END
  END cubev_ca_din0[2]
  PIN cubev_ca_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 158.480 500.000 159.080 ;
    END
  END cubev_ca_din0[30]
  PIN cubev_ca_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 161.200 500.000 161.800 ;
    END
  END cubev_ca_din0[31]
  PIN cubev_ca_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 85.040 500.000 85.640 ;
    END
  END cubev_ca_din0[3]
  PIN cubev_ca_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 87.760 500.000 88.360 ;
    END
  END cubev_ca_din0[4]
  PIN cubev_ca_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 90.480 500.000 91.080 ;
    END
  END cubev_ca_din0[5]
  PIN cubev_ca_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 93.200 500.000 93.800 ;
    END
  END cubev_ca_din0[6]
  PIN cubev_ca_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.920 500.000 96.520 ;
    END
  END cubev_ca_din0[7]
  PIN cubev_ca_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END cubev_ca_din0[8]
  PIN cubev_ca_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 101.360 500.000 101.960 ;
    END
  END cubev_ca_din0[9]
  PIN cubev_ca_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.920 500.000 164.520 ;
    END
  END cubev_ca_dout0[0]
  PIN cubev_ca_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 191.120 500.000 191.720 ;
    END
  END cubev_ca_dout0[10]
  PIN cubev_ca_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 193.840 500.000 194.440 ;
    END
  END cubev_ca_dout0[11]
  PIN cubev_ca_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 196.560 500.000 197.160 ;
    END
  END cubev_ca_dout0[12]
  PIN cubev_ca_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.280 500.000 199.880 ;
    END
  END cubev_ca_dout0[13]
  PIN cubev_ca_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 202.000 500.000 202.600 ;
    END
  END cubev_ca_dout0[14]
  PIN cubev_ca_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 204.720 500.000 205.320 ;
    END
  END cubev_ca_dout0[15]
  PIN cubev_ca_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 207.440 500.000 208.040 ;
    END
  END cubev_ca_dout0[16]
  PIN cubev_ca_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.160 500.000 210.760 ;
    END
  END cubev_ca_dout0[17]
  PIN cubev_ca_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 212.880 500.000 213.480 ;
    END
  END cubev_ca_dout0[18]
  PIN cubev_ca_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 215.600 500.000 216.200 ;
    END
  END cubev_ca_dout0[19]
  PIN cubev_ca_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END cubev_ca_dout0[1]
  PIN cubev_ca_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 218.320 500.000 218.920 ;
    END
  END cubev_ca_dout0[20]
  PIN cubev_ca_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END cubev_ca_dout0[21]
  PIN cubev_ca_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 223.760 500.000 224.360 ;
    END
  END cubev_ca_dout0[22]
  PIN cubev_ca_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 226.480 500.000 227.080 ;
    END
  END cubev_ca_dout0[23]
  PIN cubev_ca_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 229.200 500.000 229.800 ;
    END
  END cubev_ca_dout0[24]
  PIN cubev_ca_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.920 500.000 232.520 ;
    END
  END cubev_ca_dout0[25]
  PIN cubev_ca_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END cubev_ca_dout0[26]
  PIN cubev_ca_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 237.360 500.000 237.960 ;
    END
  END cubev_ca_dout0[27]
  PIN cubev_ca_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 240.080 500.000 240.680 ;
    END
  END cubev_ca_dout0[28]
  PIN cubev_ca_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 242.800 500.000 243.400 ;
    END
  END cubev_ca_dout0[29]
  PIN cubev_ca_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 169.360 500.000 169.960 ;
    END
  END cubev_ca_dout0[2]
  PIN cubev_ca_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 245.520 500.000 246.120 ;
    END
  END cubev_ca_dout0[30]
  PIN cubev_ca_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 248.240 500.000 248.840 ;
    END
  END cubev_ca_dout0[31]
  PIN cubev_ca_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 172.080 500.000 172.680 ;
    END
  END cubev_ca_dout0[3]
  PIN cubev_ca_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 174.800 500.000 175.400 ;
    END
  END cubev_ca_dout0[4]
  PIN cubev_ca_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 177.520 500.000 178.120 ;
    END
  END cubev_ca_dout0[5]
  PIN cubev_ca_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 180.240 500.000 180.840 ;
    END
  END cubev_ca_dout0[6]
  PIN cubev_ca_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 182.960 500.000 183.560 ;
    END
  END cubev_ca_dout0[7]
  PIN cubev_ca_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 185.680 500.000 186.280 ;
    END
  END cubev_ca_dout0[8]
  PIN cubev_ca_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 188.400 500.000 189.000 ;
    END
  END cubev_ca_dout0[9]
  PIN cubev_ca_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.160 500.000 278.760 ;
    END
  END cubev_ca_dout1[0]
  PIN cubev_ca_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 305.360 500.000 305.960 ;
    END
  END cubev_ca_dout1[10]
  PIN cubev_ca_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 308.080 500.000 308.680 ;
    END
  END cubev_ca_dout1[11]
  PIN cubev_ca_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 310.800 500.000 311.400 ;
    END
  END cubev_ca_dout1[12]
  PIN cubev_ca_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 313.520 500.000 314.120 ;
    END
  END cubev_ca_dout1[13]
  PIN cubev_ca_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 316.240 500.000 316.840 ;
    END
  END cubev_ca_dout1[14]
  PIN cubev_ca_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 318.960 500.000 319.560 ;
    END
  END cubev_ca_dout1[15]
  PIN cubev_ca_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 321.680 500.000 322.280 ;
    END
  END cubev_ca_dout1[16]
  PIN cubev_ca_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 324.400 500.000 325.000 ;
    END
  END cubev_ca_dout1[17]
  PIN cubev_ca_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 327.120 500.000 327.720 ;
    END
  END cubev_ca_dout1[18]
  PIN cubev_ca_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END cubev_ca_dout1[19]
  PIN cubev_ca_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 280.880 500.000 281.480 ;
    END
  END cubev_ca_dout1[1]
  PIN cubev_ca_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 332.560 500.000 333.160 ;
    END
  END cubev_ca_dout1[20]
  PIN cubev_ca_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 335.280 500.000 335.880 ;
    END
  END cubev_ca_dout1[21]
  PIN cubev_ca_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 338.000 500.000 338.600 ;
    END
  END cubev_ca_dout1[22]
  PIN cubev_ca_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.720 500.000 341.320 ;
    END
  END cubev_ca_dout1[23]
  PIN cubev_ca_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 343.440 500.000 344.040 ;
    END
  END cubev_ca_dout1[24]
  PIN cubev_ca_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 346.160 500.000 346.760 ;
    END
  END cubev_ca_dout1[25]
  PIN cubev_ca_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 348.880 500.000 349.480 ;
    END
  END cubev_ca_dout1[26]
  PIN cubev_ca_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 351.600 500.000 352.200 ;
    END
  END cubev_ca_dout1[27]
  PIN cubev_ca_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 354.320 500.000 354.920 ;
    END
  END cubev_ca_dout1[28]
  PIN cubev_ca_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END cubev_ca_dout1[29]
  PIN cubev_ca_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 283.600 500.000 284.200 ;
    END
  END cubev_ca_dout1[2]
  PIN cubev_ca_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 359.760 500.000 360.360 ;
    END
  END cubev_ca_dout1[30]
  PIN cubev_ca_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 362.480 500.000 363.080 ;
    END
  END cubev_ca_dout1[31]
  PIN cubev_ca_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 286.320 500.000 286.920 ;
    END
  END cubev_ca_dout1[3]
  PIN cubev_ca_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.040 500.000 289.640 ;
    END
  END cubev_ca_dout1[4]
  PIN cubev_ca_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 291.760 500.000 292.360 ;
    END
  END cubev_ca_dout1[5]
  PIN cubev_ca_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 294.480 500.000 295.080 ;
    END
  END cubev_ca_dout1[6]
  PIN cubev_ca_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.200 500.000 297.800 ;
    END
  END cubev_ca_dout1[7]
  PIN cubev_ca_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 299.920 500.000 300.520 ;
    END
  END cubev_ca_dout1[8]
  PIN cubev_ca_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 302.640 500.000 303.240 ;
    END
  END cubev_ca_dout1[9]
  PIN cubev_ca_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 41.520 500.000 42.120 ;
    END
  END cubev_ca_web0
  PIN cubev_ca_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END cubev_ca_wmask0[0]
  PIN cubev_ca_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 46.960 500.000 47.560 ;
    END
  END cubev_ca_wmask0[1]
  PIN cubev_ca_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 49.680 500.000 50.280 ;
    END
  END cubev_ca_wmask0[2]
  PIN cubev_ca_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 52.400 500.000 53.000 ;
    END
  END cubev_ca_wmask0[3]
  PIN cubev_phi_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 396.000 26.590 400.000 ;
    END
  END cubev_phi_addr0[0]
  PIN cubev_phi_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 396.000 29.350 400.000 ;
    END
  END cubev_phi_addr0[1]
  PIN cubev_phi_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 396.000 32.110 400.000 ;
    END
  END cubev_phi_addr0[2]
  PIN cubev_phi_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 396.000 34.870 400.000 ;
    END
  END cubev_phi_addr0[3]
  PIN cubev_phi_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 396.000 37.630 400.000 ;
    END
  END cubev_phi_addr0[4]
  PIN cubev_phi_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 396.000 40.390 400.000 ;
    END
  END cubev_phi_addr0[5]
  PIN cubev_phi_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 396.000 43.150 400.000 ;
    END
  END cubev_phi_addr0[6]
  PIN cubev_phi_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 396.000 45.910 400.000 ;
    END
  END cubev_phi_addr0[7]
  PIN cubev_phi_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 396.000 7.270 400.000 ;
    END
  END cubev_phi_clk0
  PIN cubev_phi_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 396.000 10.030 400.000 ;
    END
  END cubev_phi_csb0
  PIN cubev_phi_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END cubev_phi_din0[0]
  PIN cubev_phi_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 396.000 76.270 400.000 ;
    END
  END cubev_phi_din0[10]
  PIN cubev_phi_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 396.000 79.030 400.000 ;
    END
  END cubev_phi_din0[11]
  PIN cubev_phi_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 396.000 81.790 400.000 ;
    END
  END cubev_phi_din0[12]
  PIN cubev_phi_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 396.000 84.550 400.000 ;
    END
  END cubev_phi_din0[13]
  PIN cubev_phi_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 396.000 87.310 400.000 ;
    END
  END cubev_phi_din0[14]
  PIN cubev_phi_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 396.000 90.070 400.000 ;
    END
  END cubev_phi_din0[15]
  PIN cubev_phi_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 396.000 92.830 400.000 ;
    END
  END cubev_phi_din0[16]
  PIN cubev_phi_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 396.000 95.590 400.000 ;
    END
  END cubev_phi_din0[17]
  PIN cubev_phi_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 396.000 98.350 400.000 ;
    END
  END cubev_phi_din0[18]
  PIN cubev_phi_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 396.000 101.110 400.000 ;
    END
  END cubev_phi_din0[19]
  PIN cubev_phi_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 396.000 51.430 400.000 ;
    END
  END cubev_phi_din0[1]
  PIN cubev_phi_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 396.000 103.870 400.000 ;
    END
  END cubev_phi_din0[20]
  PIN cubev_phi_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 396.000 106.630 400.000 ;
    END
  END cubev_phi_din0[21]
  PIN cubev_phi_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 396.000 109.390 400.000 ;
    END
  END cubev_phi_din0[22]
  PIN cubev_phi_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 396.000 112.150 400.000 ;
    END
  END cubev_phi_din0[23]
  PIN cubev_phi_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 396.000 114.910 400.000 ;
    END
  END cubev_phi_din0[24]
  PIN cubev_phi_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 396.000 117.670 400.000 ;
    END
  END cubev_phi_din0[25]
  PIN cubev_phi_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 396.000 120.430 400.000 ;
    END
  END cubev_phi_din0[26]
  PIN cubev_phi_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 396.000 123.190 400.000 ;
    END
  END cubev_phi_din0[27]
  PIN cubev_phi_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 396.000 125.950 400.000 ;
    END
  END cubev_phi_din0[28]
  PIN cubev_phi_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 396.000 128.710 400.000 ;
    END
  END cubev_phi_din0[29]
  PIN cubev_phi_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 396.000 54.190 400.000 ;
    END
  END cubev_phi_din0[2]
  PIN cubev_phi_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 396.000 131.470 400.000 ;
    END
  END cubev_phi_din0[30]
  PIN cubev_phi_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 396.000 134.230 400.000 ;
    END
  END cubev_phi_din0[31]
  PIN cubev_phi_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 396.000 56.950 400.000 ;
    END
  END cubev_phi_din0[3]
  PIN cubev_phi_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END cubev_phi_din0[4]
  PIN cubev_phi_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 396.000 62.470 400.000 ;
    END
  END cubev_phi_din0[5]
  PIN cubev_phi_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 396.000 65.230 400.000 ;
    END
  END cubev_phi_din0[6]
  PIN cubev_phi_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 396.000 67.990 400.000 ;
    END
  END cubev_phi_din0[7]
  PIN cubev_phi_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 396.000 70.750 400.000 ;
    END
  END cubev_phi_din0[8]
  PIN cubev_phi_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 396.000 73.510 400.000 ;
    END
  END cubev_phi_din0[9]
  PIN cubev_phi_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 396.000 136.990 400.000 ;
    END
  END cubev_phi_dout0[0]
  PIN cubev_phi_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 396.000 164.590 400.000 ;
    END
  END cubev_phi_dout0[10]
  PIN cubev_phi_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 396.000 167.350 400.000 ;
    END
  END cubev_phi_dout0[11]
  PIN cubev_phi_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 396.000 170.110 400.000 ;
    END
  END cubev_phi_dout0[12]
  PIN cubev_phi_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 396.000 172.870 400.000 ;
    END
  END cubev_phi_dout0[13]
  PIN cubev_phi_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 396.000 175.630 400.000 ;
    END
  END cubev_phi_dout0[14]
  PIN cubev_phi_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 396.000 178.390 400.000 ;
    END
  END cubev_phi_dout0[15]
  PIN cubev_phi_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 396.000 181.150 400.000 ;
    END
  END cubev_phi_dout0[16]
  PIN cubev_phi_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 396.000 183.910 400.000 ;
    END
  END cubev_phi_dout0[17]
  PIN cubev_phi_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 396.000 186.670 400.000 ;
    END
  END cubev_phi_dout0[18]
  PIN cubev_phi_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 396.000 189.430 400.000 ;
    END
  END cubev_phi_dout0[19]
  PIN cubev_phi_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 396.000 139.750 400.000 ;
    END
  END cubev_phi_dout0[1]
  PIN cubev_phi_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 396.000 192.190 400.000 ;
    END
  END cubev_phi_dout0[20]
  PIN cubev_phi_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 396.000 194.950 400.000 ;
    END
  END cubev_phi_dout0[21]
  PIN cubev_phi_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 396.000 197.710 400.000 ;
    END
  END cubev_phi_dout0[22]
  PIN cubev_phi_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 396.000 200.470 400.000 ;
    END
  END cubev_phi_dout0[23]
  PIN cubev_phi_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 396.000 203.230 400.000 ;
    END
  END cubev_phi_dout0[24]
  PIN cubev_phi_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 396.000 205.990 400.000 ;
    END
  END cubev_phi_dout0[25]
  PIN cubev_phi_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 396.000 208.750 400.000 ;
    END
  END cubev_phi_dout0[26]
  PIN cubev_phi_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 396.000 211.510 400.000 ;
    END
  END cubev_phi_dout0[27]
  PIN cubev_phi_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 396.000 214.270 400.000 ;
    END
  END cubev_phi_dout0[28]
  PIN cubev_phi_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 396.000 217.030 400.000 ;
    END
  END cubev_phi_dout0[29]
  PIN cubev_phi_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 396.000 142.510 400.000 ;
    END
  END cubev_phi_dout0[2]
  PIN cubev_phi_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 396.000 219.790 400.000 ;
    END
  END cubev_phi_dout0[30]
  PIN cubev_phi_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 396.000 222.550 400.000 ;
    END
  END cubev_phi_dout0[31]
  PIN cubev_phi_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 396.000 145.270 400.000 ;
    END
  END cubev_phi_dout0[3]
  PIN cubev_phi_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 396.000 148.030 400.000 ;
    END
  END cubev_phi_dout0[4]
  PIN cubev_phi_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 396.000 150.790 400.000 ;
    END
  END cubev_phi_dout0[5]
  PIN cubev_phi_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 396.000 153.550 400.000 ;
    END
  END cubev_phi_dout0[6]
  PIN cubev_phi_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 396.000 156.310 400.000 ;
    END
  END cubev_phi_dout0[7]
  PIN cubev_phi_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 396.000 159.070 400.000 ;
    END
  END cubev_phi_dout0[8]
  PIN cubev_phi_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 396.000 161.830 400.000 ;
    END
  END cubev_phi_dout0[9]
  PIN cubev_phi_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 396.000 12.790 400.000 ;
    END
  END cubev_phi_web0
  PIN cubev_phi_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 396.000 15.550 400.000 ;
    END
  END cubev_phi_wmask0[0]
  PIN cubev_phi_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 396.000 18.310 400.000 ;
    END
  END cubev_phi_wmask0[1]
  PIN cubev_phi_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 396.000 21.070 400.000 ;
    END
  END cubev_phi_wmask0[2]
  PIN cubev_phi_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 396.000 23.830 400.000 ;
    END
  END cubev_phi_wmask0[3]
  PIN cubev_pli_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END cubev_pli_addr0[0]
  PIN cubev_pli_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END cubev_pli_addr0[1]
  PIN cubev_pli_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END cubev_pli_addr0[2]
  PIN cubev_pli_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END cubev_pli_addr0[3]
  PIN cubev_pli_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END cubev_pli_addr0[4]
  PIN cubev_pli_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cubev_pli_addr0[5]
  PIN cubev_pli_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END cubev_pli_addr0[6]
  PIN cubev_pli_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END cubev_pli_addr0[7]
  PIN cubev_pli_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END cubev_pli_clk0
  PIN cubev_pli_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END cubev_pli_csb0
  PIN cubev_pli_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END cubev_pli_din0[0]
  PIN cubev_pli_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END cubev_pli_din0[10]
  PIN cubev_pli_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END cubev_pli_din0[11]
  PIN cubev_pli_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END cubev_pli_din0[12]
  PIN cubev_pli_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END cubev_pli_din0[13]
  PIN cubev_pli_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END cubev_pli_din0[14]
  PIN cubev_pli_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END cubev_pli_din0[15]
  PIN cubev_pli_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END cubev_pli_din0[16]
  PIN cubev_pli_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END cubev_pli_din0[17]
  PIN cubev_pli_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END cubev_pli_din0[18]
  PIN cubev_pli_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END cubev_pli_din0[19]
  PIN cubev_pli_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END cubev_pli_din0[1]
  PIN cubev_pli_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END cubev_pli_din0[20]
  PIN cubev_pli_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END cubev_pli_din0[21]
  PIN cubev_pli_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END cubev_pli_din0[22]
  PIN cubev_pli_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END cubev_pli_din0[23]
  PIN cubev_pli_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END cubev_pli_din0[24]
  PIN cubev_pli_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END cubev_pli_din0[25]
  PIN cubev_pli_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END cubev_pli_din0[26]
  PIN cubev_pli_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END cubev_pli_din0[27]
  PIN cubev_pli_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END cubev_pli_din0[28]
  PIN cubev_pli_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END cubev_pli_din0[29]
  PIN cubev_pli_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END cubev_pli_din0[2]
  PIN cubev_pli_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END cubev_pli_din0[30]
  PIN cubev_pli_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END cubev_pli_din0[31]
  PIN cubev_pli_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END cubev_pli_din0[3]
  PIN cubev_pli_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END cubev_pli_din0[4]
  PIN cubev_pli_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END cubev_pli_din0[5]
  PIN cubev_pli_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END cubev_pli_din0[6]
  PIN cubev_pli_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END cubev_pli_din0[7]
  PIN cubev_pli_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END cubev_pli_din0[8]
  PIN cubev_pli_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END cubev_pli_din0[9]
  PIN cubev_pli_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END cubev_pli_dout0[0]
  PIN cubev_pli_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END cubev_pli_dout0[10]
  PIN cubev_pli_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END cubev_pli_dout0[11]
  PIN cubev_pli_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END cubev_pli_dout0[12]
  PIN cubev_pli_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END cubev_pli_dout0[13]
  PIN cubev_pli_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END cubev_pli_dout0[14]
  PIN cubev_pli_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END cubev_pli_dout0[15]
  PIN cubev_pli_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END cubev_pli_dout0[16]
  PIN cubev_pli_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END cubev_pli_dout0[17]
  PIN cubev_pli_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END cubev_pli_dout0[18]
  PIN cubev_pli_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END cubev_pli_dout0[19]
  PIN cubev_pli_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END cubev_pli_dout0[1]
  PIN cubev_pli_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END cubev_pli_dout0[20]
  PIN cubev_pli_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END cubev_pli_dout0[21]
  PIN cubev_pli_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END cubev_pli_dout0[22]
  PIN cubev_pli_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END cubev_pli_dout0[23]
  PIN cubev_pli_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END cubev_pli_dout0[24]
  PIN cubev_pli_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END cubev_pli_dout0[25]
  PIN cubev_pli_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END cubev_pli_dout0[26]
  PIN cubev_pli_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END cubev_pli_dout0[27]
  PIN cubev_pli_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END cubev_pli_dout0[28]
  PIN cubev_pli_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END cubev_pli_dout0[29]
  PIN cubev_pli_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END cubev_pli_dout0[2]
  PIN cubev_pli_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END cubev_pli_dout0[30]
  PIN cubev_pli_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END cubev_pli_dout0[31]
  PIN cubev_pli_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END cubev_pli_dout0[3]
  PIN cubev_pli_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END cubev_pli_dout0[4]
  PIN cubev_pli_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END cubev_pli_dout0[5]
  PIN cubev_pli_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END cubev_pli_dout0[6]
  PIN cubev_pli_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END cubev_pli_dout0[7]
  PIN cubev_pli_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END cubev_pli_dout0[8]
  PIN cubev_pli_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END cubev_pli_dout0[9]
  PIN cubev_pli_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END cubev_pli_web0
  PIN cubev_pli_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END cubev_pli_wmask0[0]
  PIN cubev_pli_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END cubev_pli_wmask0[1]
  PIN cubev_pli_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END cubev_pli_wmask0[2]
  PIN cubev_pli_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END cubev_pli_wmask0[3]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END la_oenb[9]
  PIN rstn_reg
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 396.000 493.030 400.000 ;
    END
  END rstn_reg
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 389.045 ;
      LAYER met1 ;
        RECT 5.520 5.140 494.040 391.640 ;
      LAYER met2 ;
        RECT 7.550 395.720 9.470 396.170 ;
        RECT 10.310 395.720 12.230 396.170 ;
        RECT 13.070 395.720 14.990 396.170 ;
        RECT 15.830 395.720 17.750 396.170 ;
        RECT 18.590 395.720 20.510 396.170 ;
        RECT 21.350 395.720 23.270 396.170 ;
        RECT 24.110 395.720 26.030 396.170 ;
        RECT 26.870 395.720 28.790 396.170 ;
        RECT 29.630 395.720 31.550 396.170 ;
        RECT 32.390 395.720 34.310 396.170 ;
        RECT 35.150 395.720 37.070 396.170 ;
        RECT 37.910 395.720 39.830 396.170 ;
        RECT 40.670 395.720 42.590 396.170 ;
        RECT 43.430 395.720 45.350 396.170 ;
        RECT 46.190 395.720 48.110 396.170 ;
        RECT 48.950 395.720 50.870 396.170 ;
        RECT 51.710 395.720 53.630 396.170 ;
        RECT 54.470 395.720 56.390 396.170 ;
        RECT 57.230 395.720 59.150 396.170 ;
        RECT 59.990 395.720 61.910 396.170 ;
        RECT 62.750 395.720 64.670 396.170 ;
        RECT 65.510 395.720 67.430 396.170 ;
        RECT 68.270 395.720 70.190 396.170 ;
        RECT 71.030 395.720 72.950 396.170 ;
        RECT 73.790 395.720 75.710 396.170 ;
        RECT 76.550 395.720 78.470 396.170 ;
        RECT 79.310 395.720 81.230 396.170 ;
        RECT 82.070 395.720 83.990 396.170 ;
        RECT 84.830 395.720 86.750 396.170 ;
        RECT 87.590 395.720 89.510 396.170 ;
        RECT 90.350 395.720 92.270 396.170 ;
        RECT 93.110 395.720 95.030 396.170 ;
        RECT 95.870 395.720 97.790 396.170 ;
        RECT 98.630 395.720 100.550 396.170 ;
        RECT 101.390 395.720 103.310 396.170 ;
        RECT 104.150 395.720 106.070 396.170 ;
        RECT 106.910 395.720 108.830 396.170 ;
        RECT 109.670 395.720 111.590 396.170 ;
        RECT 112.430 395.720 114.350 396.170 ;
        RECT 115.190 395.720 117.110 396.170 ;
        RECT 117.950 395.720 119.870 396.170 ;
        RECT 120.710 395.720 122.630 396.170 ;
        RECT 123.470 395.720 125.390 396.170 ;
        RECT 126.230 395.720 128.150 396.170 ;
        RECT 128.990 395.720 130.910 396.170 ;
        RECT 131.750 395.720 133.670 396.170 ;
        RECT 134.510 395.720 136.430 396.170 ;
        RECT 137.270 395.720 139.190 396.170 ;
        RECT 140.030 395.720 141.950 396.170 ;
        RECT 142.790 395.720 144.710 396.170 ;
        RECT 145.550 395.720 147.470 396.170 ;
        RECT 148.310 395.720 150.230 396.170 ;
        RECT 151.070 395.720 152.990 396.170 ;
        RECT 153.830 395.720 155.750 396.170 ;
        RECT 156.590 395.720 158.510 396.170 ;
        RECT 159.350 395.720 161.270 396.170 ;
        RECT 162.110 395.720 164.030 396.170 ;
        RECT 164.870 395.720 166.790 396.170 ;
        RECT 167.630 395.720 169.550 396.170 ;
        RECT 170.390 395.720 172.310 396.170 ;
        RECT 173.150 395.720 175.070 396.170 ;
        RECT 175.910 395.720 177.830 396.170 ;
        RECT 178.670 395.720 180.590 396.170 ;
        RECT 181.430 395.720 183.350 396.170 ;
        RECT 184.190 395.720 186.110 396.170 ;
        RECT 186.950 395.720 188.870 396.170 ;
        RECT 189.710 395.720 191.630 396.170 ;
        RECT 192.470 395.720 194.390 396.170 ;
        RECT 195.230 395.720 197.150 396.170 ;
        RECT 197.990 395.720 199.910 396.170 ;
        RECT 200.750 395.720 202.670 396.170 ;
        RECT 203.510 395.720 205.430 396.170 ;
        RECT 206.270 395.720 208.190 396.170 ;
        RECT 209.030 395.720 210.950 396.170 ;
        RECT 211.790 395.720 213.710 396.170 ;
        RECT 214.550 395.720 216.470 396.170 ;
        RECT 217.310 395.720 219.230 396.170 ;
        RECT 220.070 395.720 221.990 396.170 ;
        RECT 222.830 395.720 224.750 396.170 ;
        RECT 225.590 395.720 227.510 396.170 ;
        RECT 228.350 395.720 230.270 396.170 ;
        RECT 231.110 395.720 233.030 396.170 ;
        RECT 233.870 395.720 235.790 396.170 ;
        RECT 236.630 395.720 238.550 396.170 ;
        RECT 239.390 395.720 241.310 396.170 ;
        RECT 242.150 395.720 244.070 396.170 ;
        RECT 244.910 395.720 246.830 396.170 ;
        RECT 247.670 395.720 249.590 396.170 ;
        RECT 250.430 395.720 252.350 396.170 ;
        RECT 253.190 395.720 255.110 396.170 ;
        RECT 255.950 395.720 257.870 396.170 ;
        RECT 258.710 395.720 260.630 396.170 ;
        RECT 261.470 395.720 263.390 396.170 ;
        RECT 264.230 395.720 266.150 396.170 ;
        RECT 266.990 395.720 268.910 396.170 ;
        RECT 269.750 395.720 271.670 396.170 ;
        RECT 272.510 395.720 274.430 396.170 ;
        RECT 275.270 395.720 277.190 396.170 ;
        RECT 278.030 395.720 279.950 396.170 ;
        RECT 280.790 395.720 282.710 396.170 ;
        RECT 283.550 395.720 285.470 396.170 ;
        RECT 286.310 395.720 288.230 396.170 ;
        RECT 289.070 395.720 290.990 396.170 ;
        RECT 291.830 395.720 293.750 396.170 ;
        RECT 294.590 395.720 296.510 396.170 ;
        RECT 297.350 395.720 299.270 396.170 ;
        RECT 300.110 395.720 302.030 396.170 ;
        RECT 302.870 395.720 304.790 396.170 ;
        RECT 305.630 395.720 307.550 396.170 ;
        RECT 308.390 395.720 310.310 396.170 ;
        RECT 311.150 395.720 313.070 396.170 ;
        RECT 313.910 395.720 315.830 396.170 ;
        RECT 316.670 395.720 318.590 396.170 ;
        RECT 319.430 395.720 321.350 396.170 ;
        RECT 322.190 395.720 324.110 396.170 ;
        RECT 324.950 395.720 326.870 396.170 ;
        RECT 327.710 395.720 329.630 396.170 ;
        RECT 330.470 395.720 332.390 396.170 ;
        RECT 333.230 395.720 335.150 396.170 ;
        RECT 335.990 395.720 337.910 396.170 ;
        RECT 338.750 395.720 340.670 396.170 ;
        RECT 341.510 395.720 343.430 396.170 ;
        RECT 344.270 395.720 346.190 396.170 ;
        RECT 347.030 395.720 348.950 396.170 ;
        RECT 349.790 395.720 351.710 396.170 ;
        RECT 352.550 395.720 354.470 396.170 ;
        RECT 355.310 395.720 357.230 396.170 ;
        RECT 358.070 395.720 359.990 396.170 ;
        RECT 360.830 395.720 362.750 396.170 ;
        RECT 363.590 395.720 365.510 396.170 ;
        RECT 366.350 395.720 368.270 396.170 ;
        RECT 369.110 395.720 371.030 396.170 ;
        RECT 371.870 395.720 373.790 396.170 ;
        RECT 374.630 395.720 376.550 396.170 ;
        RECT 377.390 395.720 379.310 396.170 ;
        RECT 380.150 395.720 382.070 396.170 ;
        RECT 382.910 395.720 384.830 396.170 ;
        RECT 385.670 395.720 387.590 396.170 ;
        RECT 388.430 395.720 390.350 396.170 ;
        RECT 391.190 395.720 393.110 396.170 ;
        RECT 393.950 395.720 395.870 396.170 ;
        RECT 396.710 395.720 398.630 396.170 ;
        RECT 399.470 395.720 401.390 396.170 ;
        RECT 402.230 395.720 404.150 396.170 ;
        RECT 404.990 395.720 406.910 396.170 ;
        RECT 407.750 395.720 409.670 396.170 ;
        RECT 410.510 395.720 412.430 396.170 ;
        RECT 413.270 395.720 415.190 396.170 ;
        RECT 416.030 395.720 417.950 396.170 ;
        RECT 418.790 395.720 420.710 396.170 ;
        RECT 421.550 395.720 423.470 396.170 ;
        RECT 424.310 395.720 426.230 396.170 ;
        RECT 427.070 395.720 428.990 396.170 ;
        RECT 429.830 395.720 431.750 396.170 ;
        RECT 432.590 395.720 434.510 396.170 ;
        RECT 435.350 395.720 437.270 396.170 ;
        RECT 438.110 395.720 440.030 396.170 ;
        RECT 440.870 395.720 442.790 396.170 ;
        RECT 443.630 395.720 445.550 396.170 ;
        RECT 446.390 395.720 448.310 396.170 ;
        RECT 449.150 395.720 451.070 396.170 ;
        RECT 451.910 395.720 453.830 396.170 ;
        RECT 454.670 395.720 456.590 396.170 ;
        RECT 457.430 395.720 459.350 396.170 ;
        RECT 460.190 395.720 462.110 396.170 ;
        RECT 462.950 395.720 464.870 396.170 ;
        RECT 465.710 395.720 467.630 396.170 ;
        RECT 468.470 395.720 470.390 396.170 ;
        RECT 471.230 395.720 473.150 396.170 ;
        RECT 473.990 395.720 475.910 396.170 ;
        RECT 476.750 395.720 478.670 396.170 ;
        RECT 479.510 395.720 481.430 396.170 ;
        RECT 482.270 395.720 484.190 396.170 ;
        RECT 485.030 395.720 486.950 396.170 ;
        RECT 487.790 395.720 489.710 396.170 ;
        RECT 490.550 395.720 492.470 396.170 ;
        RECT 493.310 395.720 493.950 396.170 ;
        RECT 6.990 4.280 493.950 395.720 ;
        RECT 6.990 4.000 23.270 4.280 ;
        RECT 24.110 4.000 24.190 4.280 ;
        RECT 25.030 4.000 25.110 4.280 ;
        RECT 25.950 4.000 26.030 4.280 ;
        RECT 26.870 4.000 26.950 4.280 ;
        RECT 27.790 4.000 27.870 4.280 ;
        RECT 28.710 4.000 28.790 4.280 ;
        RECT 29.630 4.000 29.710 4.280 ;
        RECT 30.550 4.000 30.630 4.280 ;
        RECT 31.470 4.000 31.550 4.280 ;
        RECT 32.390 4.000 32.470 4.280 ;
        RECT 33.310 4.000 33.390 4.280 ;
        RECT 34.230 4.000 34.310 4.280 ;
        RECT 35.150 4.000 35.230 4.280 ;
        RECT 36.070 4.000 36.150 4.280 ;
        RECT 36.990 4.000 37.070 4.280 ;
        RECT 37.910 4.000 37.990 4.280 ;
        RECT 38.830 4.000 38.910 4.280 ;
        RECT 39.750 4.000 39.830 4.280 ;
        RECT 40.670 4.000 40.750 4.280 ;
        RECT 41.590 4.000 41.670 4.280 ;
        RECT 42.510 4.000 42.590 4.280 ;
        RECT 43.430 4.000 43.510 4.280 ;
        RECT 44.350 4.000 44.430 4.280 ;
        RECT 45.270 4.000 45.350 4.280 ;
        RECT 46.190 4.000 46.270 4.280 ;
        RECT 47.110 4.000 47.190 4.280 ;
        RECT 48.030 4.000 48.110 4.280 ;
        RECT 48.950 4.000 49.030 4.280 ;
        RECT 49.870 4.000 49.950 4.280 ;
        RECT 50.790 4.000 50.870 4.280 ;
        RECT 51.710 4.000 51.790 4.280 ;
        RECT 52.630 4.000 52.710 4.280 ;
        RECT 53.550 4.000 53.630 4.280 ;
        RECT 54.470 4.000 54.550 4.280 ;
        RECT 55.390 4.000 55.470 4.280 ;
        RECT 56.310 4.000 56.390 4.280 ;
        RECT 57.230 4.000 57.310 4.280 ;
        RECT 58.150 4.000 58.230 4.280 ;
        RECT 59.070 4.000 59.150 4.280 ;
        RECT 59.990 4.000 60.070 4.280 ;
        RECT 60.910 4.000 60.990 4.280 ;
        RECT 61.830 4.000 61.910 4.280 ;
        RECT 62.750 4.000 62.830 4.280 ;
        RECT 63.670 4.000 63.750 4.280 ;
        RECT 64.590 4.000 64.670 4.280 ;
        RECT 65.510 4.000 65.590 4.280 ;
        RECT 66.430 4.000 66.510 4.280 ;
        RECT 67.350 4.000 67.430 4.280 ;
        RECT 68.270 4.000 68.350 4.280 ;
        RECT 69.190 4.000 69.270 4.280 ;
        RECT 70.110 4.000 70.190 4.280 ;
        RECT 71.030 4.000 71.110 4.280 ;
        RECT 71.950 4.000 72.030 4.280 ;
        RECT 72.870 4.000 72.950 4.280 ;
        RECT 73.790 4.000 73.870 4.280 ;
        RECT 74.710 4.000 74.790 4.280 ;
        RECT 75.630 4.000 75.710 4.280 ;
        RECT 76.550 4.000 76.630 4.280 ;
        RECT 77.470 4.000 77.550 4.280 ;
        RECT 78.390 4.000 78.470 4.280 ;
        RECT 79.310 4.000 79.390 4.280 ;
        RECT 80.230 4.000 80.310 4.280 ;
        RECT 81.150 4.000 81.230 4.280 ;
        RECT 82.070 4.000 82.150 4.280 ;
        RECT 82.990 4.000 83.070 4.280 ;
        RECT 83.910 4.000 83.990 4.280 ;
        RECT 84.830 4.000 84.910 4.280 ;
        RECT 85.750 4.000 85.830 4.280 ;
        RECT 86.670 4.000 86.750 4.280 ;
        RECT 87.590 4.000 87.670 4.280 ;
        RECT 88.510 4.000 88.590 4.280 ;
        RECT 89.430 4.000 89.510 4.280 ;
        RECT 90.350 4.000 90.430 4.280 ;
        RECT 91.270 4.000 91.350 4.280 ;
        RECT 92.190 4.000 92.270 4.280 ;
        RECT 93.110 4.000 93.190 4.280 ;
        RECT 94.030 4.000 94.110 4.280 ;
        RECT 94.950 4.000 95.030 4.280 ;
        RECT 95.870 4.000 95.950 4.280 ;
        RECT 96.790 4.000 96.870 4.280 ;
        RECT 97.710 4.000 97.790 4.280 ;
        RECT 98.630 4.000 98.710 4.280 ;
        RECT 99.550 4.000 99.630 4.280 ;
        RECT 100.470 4.000 100.550 4.280 ;
        RECT 101.390 4.000 101.470 4.280 ;
        RECT 102.310 4.000 102.390 4.280 ;
        RECT 103.230 4.000 103.310 4.280 ;
        RECT 104.150 4.000 104.230 4.280 ;
        RECT 105.070 4.000 105.150 4.280 ;
        RECT 105.990 4.000 106.070 4.280 ;
        RECT 106.910 4.000 106.990 4.280 ;
        RECT 107.830 4.000 107.910 4.280 ;
        RECT 108.750 4.000 108.830 4.280 ;
        RECT 109.670 4.000 109.750 4.280 ;
        RECT 110.590 4.000 110.670 4.280 ;
        RECT 111.510 4.000 111.590 4.280 ;
        RECT 112.430 4.000 112.510 4.280 ;
        RECT 113.350 4.000 113.430 4.280 ;
        RECT 114.270 4.000 114.350 4.280 ;
        RECT 115.190 4.000 115.270 4.280 ;
        RECT 116.110 4.000 116.190 4.280 ;
        RECT 117.030 4.000 117.110 4.280 ;
        RECT 117.950 4.000 118.030 4.280 ;
        RECT 118.870 4.000 118.950 4.280 ;
        RECT 119.790 4.000 119.870 4.280 ;
        RECT 120.710 4.000 120.790 4.280 ;
        RECT 121.630 4.000 121.710 4.280 ;
        RECT 122.550 4.000 122.630 4.280 ;
        RECT 123.470 4.000 123.550 4.280 ;
        RECT 124.390 4.000 124.470 4.280 ;
        RECT 125.310 4.000 125.390 4.280 ;
        RECT 126.230 4.000 126.310 4.280 ;
        RECT 127.150 4.000 127.230 4.280 ;
        RECT 128.070 4.000 128.150 4.280 ;
        RECT 128.990 4.000 129.070 4.280 ;
        RECT 129.910 4.000 129.990 4.280 ;
        RECT 130.830 4.000 130.910 4.280 ;
        RECT 131.750 4.000 131.830 4.280 ;
        RECT 132.670 4.000 132.750 4.280 ;
        RECT 133.590 4.000 133.670 4.280 ;
        RECT 134.510 4.000 134.590 4.280 ;
        RECT 135.430 4.000 135.510 4.280 ;
        RECT 136.350 4.000 136.430 4.280 ;
        RECT 137.270 4.000 137.350 4.280 ;
        RECT 138.190 4.000 138.270 4.280 ;
        RECT 139.110 4.000 139.190 4.280 ;
        RECT 140.030 4.000 140.110 4.280 ;
        RECT 140.950 4.000 141.030 4.280 ;
        RECT 141.870 4.000 141.950 4.280 ;
        RECT 142.790 4.000 142.870 4.280 ;
        RECT 143.710 4.000 143.790 4.280 ;
        RECT 144.630 4.000 144.710 4.280 ;
        RECT 145.550 4.000 145.630 4.280 ;
        RECT 146.470 4.000 146.550 4.280 ;
        RECT 147.390 4.000 147.470 4.280 ;
        RECT 148.310 4.000 148.390 4.280 ;
        RECT 149.230 4.000 149.310 4.280 ;
        RECT 150.150 4.000 150.230 4.280 ;
        RECT 151.070 4.000 151.150 4.280 ;
        RECT 151.990 4.000 152.070 4.280 ;
        RECT 152.910 4.000 152.990 4.280 ;
        RECT 153.830 4.000 153.910 4.280 ;
        RECT 154.750 4.000 154.830 4.280 ;
        RECT 155.670 4.000 155.750 4.280 ;
        RECT 156.590 4.000 156.670 4.280 ;
        RECT 157.510 4.000 157.590 4.280 ;
        RECT 158.430 4.000 158.510 4.280 ;
        RECT 159.350 4.000 159.430 4.280 ;
        RECT 160.270 4.000 160.350 4.280 ;
        RECT 161.190 4.000 161.270 4.280 ;
        RECT 162.110 4.000 162.190 4.280 ;
        RECT 163.030 4.000 163.110 4.280 ;
        RECT 163.950 4.000 164.030 4.280 ;
        RECT 164.870 4.000 164.950 4.280 ;
        RECT 165.790 4.000 165.870 4.280 ;
        RECT 166.710 4.000 166.790 4.280 ;
        RECT 167.630 4.000 167.710 4.280 ;
        RECT 168.550 4.000 168.630 4.280 ;
        RECT 169.470 4.000 169.550 4.280 ;
        RECT 170.390 4.000 170.470 4.280 ;
        RECT 171.310 4.000 171.390 4.280 ;
        RECT 172.230 4.000 172.310 4.280 ;
        RECT 173.150 4.000 173.230 4.280 ;
        RECT 174.070 4.000 174.150 4.280 ;
        RECT 174.990 4.000 175.070 4.280 ;
        RECT 175.910 4.000 175.990 4.280 ;
        RECT 176.830 4.000 176.910 4.280 ;
        RECT 177.750 4.000 177.830 4.280 ;
        RECT 178.670 4.000 178.750 4.280 ;
        RECT 179.590 4.000 179.670 4.280 ;
        RECT 180.510 4.000 180.590 4.280 ;
        RECT 181.430 4.000 181.510 4.280 ;
        RECT 182.350 4.000 182.430 4.280 ;
        RECT 183.270 4.000 183.350 4.280 ;
        RECT 184.190 4.000 184.270 4.280 ;
        RECT 185.110 4.000 185.190 4.280 ;
        RECT 186.030 4.000 186.110 4.280 ;
        RECT 186.950 4.000 187.030 4.280 ;
        RECT 187.870 4.000 187.950 4.280 ;
        RECT 188.790 4.000 188.870 4.280 ;
        RECT 189.710 4.000 189.790 4.280 ;
        RECT 190.630 4.000 190.710 4.280 ;
        RECT 191.550 4.000 191.630 4.280 ;
        RECT 192.470 4.000 192.550 4.280 ;
        RECT 193.390 4.000 193.470 4.280 ;
        RECT 194.310 4.000 194.390 4.280 ;
        RECT 195.230 4.000 195.310 4.280 ;
        RECT 196.150 4.000 196.230 4.280 ;
        RECT 197.070 4.000 197.150 4.280 ;
        RECT 197.990 4.000 198.070 4.280 ;
        RECT 198.910 4.000 198.990 4.280 ;
        RECT 199.830 4.000 199.910 4.280 ;
        RECT 200.750 4.000 200.830 4.280 ;
        RECT 201.670 4.000 201.750 4.280 ;
        RECT 202.590 4.000 202.670 4.280 ;
        RECT 203.510 4.000 203.590 4.280 ;
        RECT 204.430 4.000 204.510 4.280 ;
        RECT 205.350 4.000 205.430 4.280 ;
        RECT 206.270 4.000 206.350 4.280 ;
        RECT 207.190 4.000 207.270 4.280 ;
        RECT 208.110 4.000 208.190 4.280 ;
        RECT 209.030 4.000 209.110 4.280 ;
        RECT 209.950 4.000 210.030 4.280 ;
        RECT 210.870 4.000 210.950 4.280 ;
        RECT 211.790 4.000 211.870 4.280 ;
        RECT 212.710 4.000 212.790 4.280 ;
        RECT 213.630 4.000 213.710 4.280 ;
        RECT 214.550 4.000 214.630 4.280 ;
        RECT 215.470 4.000 215.550 4.280 ;
        RECT 216.390 4.000 216.470 4.280 ;
        RECT 217.310 4.000 217.390 4.280 ;
        RECT 218.230 4.000 218.310 4.280 ;
        RECT 219.150 4.000 219.230 4.280 ;
        RECT 220.070 4.000 220.150 4.280 ;
        RECT 220.990 4.000 221.070 4.280 ;
        RECT 221.910 4.000 221.990 4.280 ;
        RECT 222.830 4.000 222.910 4.280 ;
        RECT 223.750 4.000 223.830 4.280 ;
        RECT 224.670 4.000 224.750 4.280 ;
        RECT 225.590 4.000 225.670 4.280 ;
        RECT 226.510 4.000 226.590 4.280 ;
        RECT 227.430 4.000 227.510 4.280 ;
        RECT 228.350 4.000 228.430 4.280 ;
        RECT 229.270 4.000 229.350 4.280 ;
        RECT 230.190 4.000 230.270 4.280 ;
        RECT 231.110 4.000 231.190 4.280 ;
        RECT 232.030 4.000 232.110 4.280 ;
        RECT 232.950 4.000 233.030 4.280 ;
        RECT 233.870 4.000 233.950 4.280 ;
        RECT 234.790 4.000 234.870 4.280 ;
        RECT 235.710 4.000 235.790 4.280 ;
        RECT 236.630 4.000 236.710 4.280 ;
        RECT 237.550 4.000 237.630 4.280 ;
        RECT 238.470 4.000 238.550 4.280 ;
        RECT 239.390 4.000 239.470 4.280 ;
        RECT 240.310 4.000 240.390 4.280 ;
        RECT 241.230 4.000 241.310 4.280 ;
        RECT 242.150 4.000 242.230 4.280 ;
        RECT 243.070 4.000 243.150 4.280 ;
        RECT 243.990 4.000 244.070 4.280 ;
        RECT 244.910 4.000 244.990 4.280 ;
        RECT 245.830 4.000 245.910 4.280 ;
        RECT 246.750 4.000 246.830 4.280 ;
        RECT 247.670 4.000 247.750 4.280 ;
        RECT 248.590 4.000 248.670 4.280 ;
        RECT 249.510 4.000 249.590 4.280 ;
        RECT 250.430 4.000 250.510 4.280 ;
        RECT 251.350 4.000 251.430 4.280 ;
        RECT 252.270 4.000 252.350 4.280 ;
        RECT 253.190 4.000 253.270 4.280 ;
        RECT 254.110 4.000 254.190 4.280 ;
        RECT 255.030 4.000 255.110 4.280 ;
        RECT 255.950 4.000 256.030 4.280 ;
        RECT 256.870 4.000 256.950 4.280 ;
        RECT 257.790 4.000 257.870 4.280 ;
        RECT 258.710 4.000 258.790 4.280 ;
        RECT 259.630 4.000 259.710 4.280 ;
        RECT 260.550 4.000 260.630 4.280 ;
        RECT 261.470 4.000 261.550 4.280 ;
        RECT 262.390 4.000 262.470 4.280 ;
        RECT 263.310 4.000 263.390 4.280 ;
        RECT 264.230 4.000 264.310 4.280 ;
        RECT 265.150 4.000 265.230 4.280 ;
        RECT 266.070 4.000 266.150 4.280 ;
        RECT 266.990 4.000 267.070 4.280 ;
        RECT 267.910 4.000 267.990 4.280 ;
        RECT 268.830 4.000 268.910 4.280 ;
        RECT 269.750 4.000 269.830 4.280 ;
        RECT 270.670 4.000 270.750 4.280 ;
        RECT 271.590 4.000 271.670 4.280 ;
        RECT 272.510 4.000 272.590 4.280 ;
        RECT 273.430 4.000 273.510 4.280 ;
        RECT 274.350 4.000 274.430 4.280 ;
        RECT 275.270 4.000 275.350 4.280 ;
        RECT 276.190 4.000 276.270 4.280 ;
        RECT 277.110 4.000 277.190 4.280 ;
        RECT 278.030 4.000 278.110 4.280 ;
        RECT 278.950 4.000 279.030 4.280 ;
        RECT 279.870 4.000 279.950 4.280 ;
        RECT 280.790 4.000 280.870 4.280 ;
        RECT 281.710 4.000 281.790 4.280 ;
        RECT 282.630 4.000 282.710 4.280 ;
        RECT 283.550 4.000 283.630 4.280 ;
        RECT 284.470 4.000 284.550 4.280 ;
        RECT 285.390 4.000 285.470 4.280 ;
        RECT 286.310 4.000 286.390 4.280 ;
        RECT 287.230 4.000 287.310 4.280 ;
        RECT 288.150 4.000 288.230 4.280 ;
        RECT 289.070 4.000 289.150 4.280 ;
        RECT 289.990 4.000 290.070 4.280 ;
        RECT 290.910 4.000 290.990 4.280 ;
        RECT 291.830 4.000 291.910 4.280 ;
        RECT 292.750 4.000 292.830 4.280 ;
        RECT 293.670 4.000 293.750 4.280 ;
        RECT 294.590 4.000 294.670 4.280 ;
        RECT 295.510 4.000 295.590 4.280 ;
        RECT 296.430 4.000 296.510 4.280 ;
        RECT 297.350 4.000 297.430 4.280 ;
        RECT 298.270 4.000 298.350 4.280 ;
        RECT 299.190 4.000 299.270 4.280 ;
        RECT 300.110 4.000 300.190 4.280 ;
        RECT 301.030 4.000 301.110 4.280 ;
        RECT 301.950 4.000 302.030 4.280 ;
        RECT 302.870 4.000 302.950 4.280 ;
        RECT 303.790 4.000 303.870 4.280 ;
        RECT 304.710 4.000 304.790 4.280 ;
        RECT 305.630 4.000 305.710 4.280 ;
        RECT 306.550 4.000 306.630 4.280 ;
        RECT 307.470 4.000 307.550 4.280 ;
        RECT 308.390 4.000 308.470 4.280 ;
        RECT 309.310 4.000 309.390 4.280 ;
        RECT 310.230 4.000 310.310 4.280 ;
        RECT 311.150 4.000 311.230 4.280 ;
        RECT 312.070 4.000 312.150 4.280 ;
        RECT 312.990 4.000 313.070 4.280 ;
        RECT 313.910 4.000 313.990 4.280 ;
        RECT 314.830 4.000 314.910 4.280 ;
        RECT 315.750 4.000 315.830 4.280 ;
        RECT 316.670 4.000 316.750 4.280 ;
        RECT 317.590 4.000 317.670 4.280 ;
        RECT 318.510 4.000 318.590 4.280 ;
        RECT 319.430 4.000 319.510 4.280 ;
        RECT 320.350 4.000 320.430 4.280 ;
        RECT 321.270 4.000 321.350 4.280 ;
        RECT 322.190 4.000 322.270 4.280 ;
        RECT 323.110 4.000 323.190 4.280 ;
        RECT 324.030 4.000 324.110 4.280 ;
        RECT 324.950 4.000 325.030 4.280 ;
        RECT 325.870 4.000 325.950 4.280 ;
        RECT 326.790 4.000 326.870 4.280 ;
        RECT 327.710 4.000 327.790 4.280 ;
        RECT 328.630 4.000 328.710 4.280 ;
        RECT 329.550 4.000 329.630 4.280 ;
        RECT 330.470 4.000 330.550 4.280 ;
        RECT 331.390 4.000 331.470 4.280 ;
        RECT 332.310 4.000 332.390 4.280 ;
        RECT 333.230 4.000 333.310 4.280 ;
        RECT 334.150 4.000 334.230 4.280 ;
        RECT 335.070 4.000 335.150 4.280 ;
        RECT 335.990 4.000 336.070 4.280 ;
        RECT 336.910 4.000 336.990 4.280 ;
        RECT 337.830 4.000 337.910 4.280 ;
        RECT 338.750 4.000 338.830 4.280 ;
        RECT 339.670 4.000 339.750 4.280 ;
        RECT 340.590 4.000 340.670 4.280 ;
        RECT 341.510 4.000 341.590 4.280 ;
        RECT 342.430 4.000 342.510 4.280 ;
        RECT 343.350 4.000 343.430 4.280 ;
        RECT 344.270 4.000 344.350 4.280 ;
        RECT 345.190 4.000 345.270 4.280 ;
        RECT 346.110 4.000 346.190 4.280 ;
        RECT 347.030 4.000 347.110 4.280 ;
        RECT 347.950 4.000 348.030 4.280 ;
        RECT 348.870 4.000 348.950 4.280 ;
        RECT 349.790 4.000 349.870 4.280 ;
        RECT 350.710 4.000 350.790 4.280 ;
        RECT 351.630 4.000 351.710 4.280 ;
        RECT 352.550 4.000 352.630 4.280 ;
        RECT 353.470 4.000 353.550 4.280 ;
        RECT 354.390 4.000 354.470 4.280 ;
        RECT 355.310 4.000 355.390 4.280 ;
        RECT 356.230 4.000 356.310 4.280 ;
        RECT 357.150 4.000 357.230 4.280 ;
        RECT 358.070 4.000 358.150 4.280 ;
        RECT 358.990 4.000 359.070 4.280 ;
        RECT 359.910 4.000 359.990 4.280 ;
        RECT 360.830 4.000 360.910 4.280 ;
        RECT 361.750 4.000 361.830 4.280 ;
        RECT 362.670 4.000 362.750 4.280 ;
        RECT 363.590 4.000 363.670 4.280 ;
        RECT 364.510 4.000 364.590 4.280 ;
        RECT 365.430 4.000 365.510 4.280 ;
        RECT 366.350 4.000 366.430 4.280 ;
        RECT 367.270 4.000 367.350 4.280 ;
        RECT 368.190 4.000 368.270 4.280 ;
        RECT 369.110 4.000 369.190 4.280 ;
        RECT 370.030 4.000 370.110 4.280 ;
        RECT 370.950 4.000 371.030 4.280 ;
        RECT 371.870 4.000 371.950 4.280 ;
        RECT 372.790 4.000 372.870 4.280 ;
        RECT 373.710 4.000 373.790 4.280 ;
        RECT 374.630 4.000 374.710 4.280 ;
        RECT 375.550 4.000 375.630 4.280 ;
        RECT 376.470 4.000 376.550 4.280 ;
        RECT 377.390 4.000 377.470 4.280 ;
        RECT 378.310 4.000 378.390 4.280 ;
        RECT 379.230 4.000 379.310 4.280 ;
        RECT 380.150 4.000 380.230 4.280 ;
        RECT 381.070 4.000 381.150 4.280 ;
        RECT 381.990 4.000 382.070 4.280 ;
        RECT 382.910 4.000 382.990 4.280 ;
        RECT 383.830 4.000 383.910 4.280 ;
        RECT 384.750 4.000 384.830 4.280 ;
        RECT 385.670 4.000 385.750 4.280 ;
        RECT 386.590 4.000 386.670 4.280 ;
        RECT 387.510 4.000 387.590 4.280 ;
        RECT 388.430 4.000 388.510 4.280 ;
        RECT 389.350 4.000 389.430 4.280 ;
        RECT 390.270 4.000 390.350 4.280 ;
        RECT 391.190 4.000 391.270 4.280 ;
        RECT 392.110 4.000 392.190 4.280 ;
        RECT 393.030 4.000 393.110 4.280 ;
        RECT 393.950 4.000 394.030 4.280 ;
        RECT 394.870 4.000 394.950 4.280 ;
        RECT 395.790 4.000 395.870 4.280 ;
        RECT 396.710 4.000 396.790 4.280 ;
        RECT 397.630 4.000 397.710 4.280 ;
        RECT 398.550 4.000 398.630 4.280 ;
        RECT 399.470 4.000 399.550 4.280 ;
        RECT 400.390 4.000 400.470 4.280 ;
        RECT 401.310 4.000 401.390 4.280 ;
        RECT 402.230 4.000 402.310 4.280 ;
        RECT 403.150 4.000 403.230 4.280 ;
        RECT 404.070 4.000 404.150 4.280 ;
        RECT 404.990 4.000 405.070 4.280 ;
        RECT 405.910 4.000 405.990 4.280 ;
        RECT 406.830 4.000 406.910 4.280 ;
        RECT 407.750 4.000 407.830 4.280 ;
        RECT 408.670 4.000 408.750 4.280 ;
        RECT 409.590 4.000 409.670 4.280 ;
        RECT 410.510 4.000 410.590 4.280 ;
        RECT 411.430 4.000 411.510 4.280 ;
        RECT 412.350 4.000 412.430 4.280 ;
        RECT 413.270 4.000 413.350 4.280 ;
        RECT 414.190 4.000 414.270 4.280 ;
        RECT 415.110 4.000 415.190 4.280 ;
        RECT 416.030 4.000 416.110 4.280 ;
        RECT 416.950 4.000 417.030 4.280 ;
        RECT 417.870 4.000 417.950 4.280 ;
        RECT 418.790 4.000 418.870 4.280 ;
        RECT 419.710 4.000 419.790 4.280 ;
        RECT 420.630 4.000 420.710 4.280 ;
        RECT 421.550 4.000 421.630 4.280 ;
        RECT 422.470 4.000 422.550 4.280 ;
        RECT 423.390 4.000 423.470 4.280 ;
        RECT 424.310 4.000 424.390 4.280 ;
        RECT 425.230 4.000 425.310 4.280 ;
        RECT 426.150 4.000 426.230 4.280 ;
        RECT 427.070 4.000 427.150 4.280 ;
        RECT 427.990 4.000 428.070 4.280 ;
        RECT 428.910 4.000 428.990 4.280 ;
        RECT 429.830 4.000 429.910 4.280 ;
        RECT 430.750 4.000 430.830 4.280 ;
        RECT 431.670 4.000 431.750 4.280 ;
        RECT 432.590 4.000 432.670 4.280 ;
        RECT 433.510 4.000 433.590 4.280 ;
        RECT 434.430 4.000 434.510 4.280 ;
        RECT 435.350 4.000 435.430 4.280 ;
        RECT 436.270 4.000 436.350 4.280 ;
        RECT 437.190 4.000 437.270 4.280 ;
        RECT 438.110 4.000 438.190 4.280 ;
        RECT 439.030 4.000 439.110 4.280 ;
        RECT 439.950 4.000 440.030 4.280 ;
        RECT 440.870 4.000 440.950 4.280 ;
        RECT 441.790 4.000 441.870 4.280 ;
        RECT 442.710 4.000 442.790 4.280 ;
        RECT 443.630 4.000 443.710 4.280 ;
        RECT 444.550 4.000 444.630 4.280 ;
        RECT 445.470 4.000 445.550 4.280 ;
        RECT 446.390 4.000 446.470 4.280 ;
        RECT 447.310 4.000 447.390 4.280 ;
        RECT 448.230 4.000 448.310 4.280 ;
        RECT 449.150 4.000 449.230 4.280 ;
        RECT 450.070 4.000 450.150 4.280 ;
        RECT 450.990 4.000 451.070 4.280 ;
        RECT 451.910 4.000 451.990 4.280 ;
        RECT 452.830 4.000 452.910 4.280 ;
        RECT 453.750 4.000 453.830 4.280 ;
        RECT 454.670 4.000 454.750 4.280 ;
        RECT 455.590 4.000 455.670 4.280 ;
        RECT 456.510 4.000 456.590 4.280 ;
        RECT 457.430 4.000 457.510 4.280 ;
        RECT 458.350 4.000 458.430 4.280 ;
        RECT 459.270 4.000 459.350 4.280 ;
        RECT 460.190 4.000 460.270 4.280 ;
        RECT 461.110 4.000 461.190 4.280 ;
        RECT 462.030 4.000 462.110 4.280 ;
        RECT 462.950 4.000 463.030 4.280 ;
        RECT 463.870 4.000 463.950 4.280 ;
        RECT 464.790 4.000 464.870 4.280 ;
        RECT 465.710 4.000 465.790 4.280 ;
        RECT 466.630 4.000 466.710 4.280 ;
        RECT 467.550 4.000 467.630 4.280 ;
        RECT 468.470 4.000 468.550 4.280 ;
        RECT 469.390 4.000 469.470 4.280 ;
        RECT 470.310 4.000 470.390 4.280 ;
        RECT 471.230 4.000 471.310 4.280 ;
        RECT 472.150 4.000 472.230 4.280 ;
        RECT 473.070 4.000 473.150 4.280 ;
        RECT 473.990 4.000 474.070 4.280 ;
        RECT 474.910 4.000 474.990 4.280 ;
        RECT 475.830 4.000 475.910 4.280 ;
        RECT 476.750 4.000 493.950 4.280 ;
      LAYER met3 ;
        RECT 4.000 385.920 496.000 389.125 ;
        RECT 4.400 384.520 496.000 385.920 ;
        RECT 4.000 381.160 496.000 384.520 ;
        RECT 4.400 379.760 496.000 381.160 ;
        RECT 4.000 376.400 496.000 379.760 ;
        RECT 4.400 375.000 496.000 376.400 ;
        RECT 4.000 371.640 496.000 375.000 ;
        RECT 4.400 370.240 496.000 371.640 ;
        RECT 4.000 366.880 496.000 370.240 ;
        RECT 4.400 365.480 496.000 366.880 ;
        RECT 4.000 363.480 496.000 365.480 ;
        RECT 4.000 362.120 495.600 363.480 ;
        RECT 4.400 362.080 495.600 362.120 ;
        RECT 4.400 360.760 496.000 362.080 ;
        RECT 4.400 360.720 495.600 360.760 ;
        RECT 4.000 359.360 495.600 360.720 ;
        RECT 4.000 358.040 496.000 359.360 ;
        RECT 4.000 357.360 495.600 358.040 ;
        RECT 4.400 356.640 495.600 357.360 ;
        RECT 4.400 355.960 496.000 356.640 ;
        RECT 4.000 355.320 496.000 355.960 ;
        RECT 4.000 353.920 495.600 355.320 ;
        RECT 4.000 352.600 496.000 353.920 ;
        RECT 4.400 351.200 495.600 352.600 ;
        RECT 4.000 349.880 496.000 351.200 ;
        RECT 4.000 348.480 495.600 349.880 ;
        RECT 4.000 347.840 496.000 348.480 ;
        RECT 4.400 347.160 496.000 347.840 ;
        RECT 4.400 346.440 495.600 347.160 ;
        RECT 4.000 345.760 495.600 346.440 ;
        RECT 4.000 344.440 496.000 345.760 ;
        RECT 4.000 343.080 495.600 344.440 ;
        RECT 4.400 343.040 495.600 343.080 ;
        RECT 4.400 341.720 496.000 343.040 ;
        RECT 4.400 341.680 495.600 341.720 ;
        RECT 4.000 340.320 495.600 341.680 ;
        RECT 4.000 339.000 496.000 340.320 ;
        RECT 4.000 338.320 495.600 339.000 ;
        RECT 4.400 337.600 495.600 338.320 ;
        RECT 4.400 336.920 496.000 337.600 ;
        RECT 4.000 336.280 496.000 336.920 ;
        RECT 4.000 334.880 495.600 336.280 ;
        RECT 4.000 333.560 496.000 334.880 ;
        RECT 4.400 332.160 495.600 333.560 ;
        RECT 4.000 330.840 496.000 332.160 ;
        RECT 4.000 329.440 495.600 330.840 ;
        RECT 4.000 328.800 496.000 329.440 ;
        RECT 4.400 328.120 496.000 328.800 ;
        RECT 4.400 327.400 495.600 328.120 ;
        RECT 4.000 326.720 495.600 327.400 ;
        RECT 4.000 325.400 496.000 326.720 ;
        RECT 4.000 324.040 495.600 325.400 ;
        RECT 4.400 324.000 495.600 324.040 ;
        RECT 4.400 322.680 496.000 324.000 ;
        RECT 4.400 322.640 495.600 322.680 ;
        RECT 4.000 321.280 495.600 322.640 ;
        RECT 4.000 319.960 496.000 321.280 ;
        RECT 4.000 319.280 495.600 319.960 ;
        RECT 4.400 318.560 495.600 319.280 ;
        RECT 4.400 317.880 496.000 318.560 ;
        RECT 4.000 317.240 496.000 317.880 ;
        RECT 4.000 315.840 495.600 317.240 ;
        RECT 4.000 314.520 496.000 315.840 ;
        RECT 4.400 313.120 495.600 314.520 ;
        RECT 4.000 311.800 496.000 313.120 ;
        RECT 4.000 310.400 495.600 311.800 ;
        RECT 4.000 309.760 496.000 310.400 ;
        RECT 4.400 309.080 496.000 309.760 ;
        RECT 4.400 308.360 495.600 309.080 ;
        RECT 4.000 307.680 495.600 308.360 ;
        RECT 4.000 306.360 496.000 307.680 ;
        RECT 4.000 305.000 495.600 306.360 ;
        RECT 4.400 304.960 495.600 305.000 ;
        RECT 4.400 303.640 496.000 304.960 ;
        RECT 4.400 303.600 495.600 303.640 ;
        RECT 4.000 302.240 495.600 303.600 ;
        RECT 4.000 300.920 496.000 302.240 ;
        RECT 4.000 300.240 495.600 300.920 ;
        RECT 4.400 299.520 495.600 300.240 ;
        RECT 4.400 298.840 496.000 299.520 ;
        RECT 4.000 298.200 496.000 298.840 ;
        RECT 4.000 296.800 495.600 298.200 ;
        RECT 4.000 295.480 496.000 296.800 ;
        RECT 4.400 294.080 495.600 295.480 ;
        RECT 4.000 292.760 496.000 294.080 ;
        RECT 4.000 291.360 495.600 292.760 ;
        RECT 4.000 290.720 496.000 291.360 ;
        RECT 4.400 290.040 496.000 290.720 ;
        RECT 4.400 289.320 495.600 290.040 ;
        RECT 4.000 288.640 495.600 289.320 ;
        RECT 4.000 287.320 496.000 288.640 ;
        RECT 4.000 285.960 495.600 287.320 ;
        RECT 4.400 285.920 495.600 285.960 ;
        RECT 4.400 284.600 496.000 285.920 ;
        RECT 4.400 284.560 495.600 284.600 ;
        RECT 4.000 283.200 495.600 284.560 ;
        RECT 4.000 281.880 496.000 283.200 ;
        RECT 4.000 281.200 495.600 281.880 ;
        RECT 4.400 280.480 495.600 281.200 ;
        RECT 4.400 279.800 496.000 280.480 ;
        RECT 4.000 279.160 496.000 279.800 ;
        RECT 4.000 277.760 495.600 279.160 ;
        RECT 4.000 276.440 496.000 277.760 ;
        RECT 4.400 275.040 495.600 276.440 ;
        RECT 4.000 273.720 496.000 275.040 ;
        RECT 4.000 272.320 495.600 273.720 ;
        RECT 4.000 271.680 496.000 272.320 ;
        RECT 4.400 271.000 496.000 271.680 ;
        RECT 4.400 270.280 495.600 271.000 ;
        RECT 4.000 269.600 495.600 270.280 ;
        RECT 4.000 268.280 496.000 269.600 ;
        RECT 4.000 266.920 495.600 268.280 ;
        RECT 4.400 266.880 495.600 266.920 ;
        RECT 4.400 265.560 496.000 266.880 ;
        RECT 4.400 265.520 495.600 265.560 ;
        RECT 4.000 264.160 495.600 265.520 ;
        RECT 4.000 262.840 496.000 264.160 ;
        RECT 4.000 262.160 495.600 262.840 ;
        RECT 4.400 261.440 495.600 262.160 ;
        RECT 4.400 260.760 496.000 261.440 ;
        RECT 4.000 260.120 496.000 260.760 ;
        RECT 4.000 258.720 495.600 260.120 ;
        RECT 4.000 257.400 496.000 258.720 ;
        RECT 4.400 256.000 495.600 257.400 ;
        RECT 4.000 254.680 496.000 256.000 ;
        RECT 4.000 253.280 495.600 254.680 ;
        RECT 4.000 252.640 496.000 253.280 ;
        RECT 4.400 251.960 496.000 252.640 ;
        RECT 4.400 251.240 495.600 251.960 ;
        RECT 4.000 250.560 495.600 251.240 ;
        RECT 4.000 249.240 496.000 250.560 ;
        RECT 4.000 247.880 495.600 249.240 ;
        RECT 4.400 247.840 495.600 247.880 ;
        RECT 4.400 246.520 496.000 247.840 ;
        RECT 4.400 246.480 495.600 246.520 ;
        RECT 4.000 245.120 495.600 246.480 ;
        RECT 4.000 243.800 496.000 245.120 ;
        RECT 4.000 243.120 495.600 243.800 ;
        RECT 4.400 242.400 495.600 243.120 ;
        RECT 4.400 241.720 496.000 242.400 ;
        RECT 4.000 241.080 496.000 241.720 ;
        RECT 4.000 239.680 495.600 241.080 ;
        RECT 4.000 238.360 496.000 239.680 ;
        RECT 4.400 236.960 495.600 238.360 ;
        RECT 4.000 235.640 496.000 236.960 ;
        RECT 4.000 234.240 495.600 235.640 ;
        RECT 4.000 233.600 496.000 234.240 ;
        RECT 4.400 232.920 496.000 233.600 ;
        RECT 4.400 232.200 495.600 232.920 ;
        RECT 4.000 231.520 495.600 232.200 ;
        RECT 4.000 230.200 496.000 231.520 ;
        RECT 4.000 228.840 495.600 230.200 ;
        RECT 4.400 228.800 495.600 228.840 ;
        RECT 4.400 227.480 496.000 228.800 ;
        RECT 4.400 227.440 495.600 227.480 ;
        RECT 4.000 226.080 495.600 227.440 ;
        RECT 4.000 224.760 496.000 226.080 ;
        RECT 4.000 224.080 495.600 224.760 ;
        RECT 4.400 223.360 495.600 224.080 ;
        RECT 4.400 222.680 496.000 223.360 ;
        RECT 4.000 222.040 496.000 222.680 ;
        RECT 4.000 220.640 495.600 222.040 ;
        RECT 4.000 219.320 496.000 220.640 ;
        RECT 4.400 217.920 495.600 219.320 ;
        RECT 4.000 216.600 496.000 217.920 ;
        RECT 4.000 215.200 495.600 216.600 ;
        RECT 4.000 214.560 496.000 215.200 ;
        RECT 4.400 213.880 496.000 214.560 ;
        RECT 4.400 213.160 495.600 213.880 ;
        RECT 4.000 212.480 495.600 213.160 ;
        RECT 4.000 211.160 496.000 212.480 ;
        RECT 4.000 209.800 495.600 211.160 ;
        RECT 4.400 209.760 495.600 209.800 ;
        RECT 4.400 208.440 496.000 209.760 ;
        RECT 4.400 208.400 495.600 208.440 ;
        RECT 4.000 207.040 495.600 208.400 ;
        RECT 4.000 205.720 496.000 207.040 ;
        RECT 4.000 205.040 495.600 205.720 ;
        RECT 4.400 204.320 495.600 205.040 ;
        RECT 4.400 203.640 496.000 204.320 ;
        RECT 4.000 203.000 496.000 203.640 ;
        RECT 4.000 201.600 495.600 203.000 ;
        RECT 4.000 200.280 496.000 201.600 ;
        RECT 4.400 198.880 495.600 200.280 ;
        RECT 4.000 197.560 496.000 198.880 ;
        RECT 4.000 196.160 495.600 197.560 ;
        RECT 4.000 195.520 496.000 196.160 ;
        RECT 4.400 194.840 496.000 195.520 ;
        RECT 4.400 194.120 495.600 194.840 ;
        RECT 4.000 193.440 495.600 194.120 ;
        RECT 4.000 192.120 496.000 193.440 ;
        RECT 4.000 190.760 495.600 192.120 ;
        RECT 4.400 190.720 495.600 190.760 ;
        RECT 4.400 189.400 496.000 190.720 ;
        RECT 4.400 189.360 495.600 189.400 ;
        RECT 4.000 188.000 495.600 189.360 ;
        RECT 4.000 186.680 496.000 188.000 ;
        RECT 4.000 186.000 495.600 186.680 ;
        RECT 4.400 185.280 495.600 186.000 ;
        RECT 4.400 184.600 496.000 185.280 ;
        RECT 4.000 183.960 496.000 184.600 ;
        RECT 4.000 182.560 495.600 183.960 ;
        RECT 4.000 181.240 496.000 182.560 ;
        RECT 4.400 179.840 495.600 181.240 ;
        RECT 4.000 178.520 496.000 179.840 ;
        RECT 4.000 177.120 495.600 178.520 ;
        RECT 4.000 176.480 496.000 177.120 ;
        RECT 4.400 175.800 496.000 176.480 ;
        RECT 4.400 175.080 495.600 175.800 ;
        RECT 4.000 174.400 495.600 175.080 ;
        RECT 4.000 173.080 496.000 174.400 ;
        RECT 4.000 171.720 495.600 173.080 ;
        RECT 4.400 171.680 495.600 171.720 ;
        RECT 4.400 170.360 496.000 171.680 ;
        RECT 4.400 170.320 495.600 170.360 ;
        RECT 4.000 168.960 495.600 170.320 ;
        RECT 4.000 167.640 496.000 168.960 ;
        RECT 4.000 166.960 495.600 167.640 ;
        RECT 4.400 166.240 495.600 166.960 ;
        RECT 4.400 165.560 496.000 166.240 ;
        RECT 4.000 164.920 496.000 165.560 ;
        RECT 4.000 163.520 495.600 164.920 ;
        RECT 4.000 162.200 496.000 163.520 ;
        RECT 4.400 160.800 495.600 162.200 ;
        RECT 4.000 159.480 496.000 160.800 ;
        RECT 4.000 158.080 495.600 159.480 ;
        RECT 4.000 157.440 496.000 158.080 ;
        RECT 4.400 156.760 496.000 157.440 ;
        RECT 4.400 156.040 495.600 156.760 ;
        RECT 4.000 155.360 495.600 156.040 ;
        RECT 4.000 154.040 496.000 155.360 ;
        RECT 4.000 152.680 495.600 154.040 ;
        RECT 4.400 152.640 495.600 152.680 ;
        RECT 4.400 151.320 496.000 152.640 ;
        RECT 4.400 151.280 495.600 151.320 ;
        RECT 4.000 149.920 495.600 151.280 ;
        RECT 4.000 148.600 496.000 149.920 ;
        RECT 4.000 147.920 495.600 148.600 ;
        RECT 4.400 147.200 495.600 147.920 ;
        RECT 4.400 146.520 496.000 147.200 ;
        RECT 4.000 145.880 496.000 146.520 ;
        RECT 4.000 144.480 495.600 145.880 ;
        RECT 4.000 143.160 496.000 144.480 ;
        RECT 4.400 141.760 495.600 143.160 ;
        RECT 4.000 140.440 496.000 141.760 ;
        RECT 4.000 139.040 495.600 140.440 ;
        RECT 4.000 138.400 496.000 139.040 ;
        RECT 4.400 137.720 496.000 138.400 ;
        RECT 4.400 137.000 495.600 137.720 ;
        RECT 4.000 136.320 495.600 137.000 ;
        RECT 4.000 135.000 496.000 136.320 ;
        RECT 4.000 133.640 495.600 135.000 ;
        RECT 4.400 133.600 495.600 133.640 ;
        RECT 4.400 132.280 496.000 133.600 ;
        RECT 4.400 132.240 495.600 132.280 ;
        RECT 4.000 130.880 495.600 132.240 ;
        RECT 4.000 129.560 496.000 130.880 ;
        RECT 4.000 128.880 495.600 129.560 ;
        RECT 4.400 128.160 495.600 128.880 ;
        RECT 4.400 127.480 496.000 128.160 ;
        RECT 4.000 126.840 496.000 127.480 ;
        RECT 4.000 125.440 495.600 126.840 ;
        RECT 4.000 124.120 496.000 125.440 ;
        RECT 4.400 122.720 495.600 124.120 ;
        RECT 4.000 121.400 496.000 122.720 ;
        RECT 4.000 120.000 495.600 121.400 ;
        RECT 4.000 119.360 496.000 120.000 ;
        RECT 4.400 118.680 496.000 119.360 ;
        RECT 4.400 117.960 495.600 118.680 ;
        RECT 4.000 117.280 495.600 117.960 ;
        RECT 4.000 115.960 496.000 117.280 ;
        RECT 4.000 114.600 495.600 115.960 ;
        RECT 4.400 114.560 495.600 114.600 ;
        RECT 4.400 113.240 496.000 114.560 ;
        RECT 4.400 113.200 495.600 113.240 ;
        RECT 4.000 111.840 495.600 113.200 ;
        RECT 4.000 110.520 496.000 111.840 ;
        RECT 4.000 109.840 495.600 110.520 ;
        RECT 4.400 109.120 495.600 109.840 ;
        RECT 4.400 108.440 496.000 109.120 ;
        RECT 4.000 107.800 496.000 108.440 ;
        RECT 4.000 106.400 495.600 107.800 ;
        RECT 4.000 105.080 496.000 106.400 ;
        RECT 4.400 103.680 495.600 105.080 ;
        RECT 4.000 102.360 496.000 103.680 ;
        RECT 4.000 100.960 495.600 102.360 ;
        RECT 4.000 100.320 496.000 100.960 ;
        RECT 4.400 99.640 496.000 100.320 ;
        RECT 4.400 98.920 495.600 99.640 ;
        RECT 4.000 98.240 495.600 98.920 ;
        RECT 4.000 96.920 496.000 98.240 ;
        RECT 4.000 95.560 495.600 96.920 ;
        RECT 4.400 95.520 495.600 95.560 ;
        RECT 4.400 94.200 496.000 95.520 ;
        RECT 4.400 94.160 495.600 94.200 ;
        RECT 4.000 92.800 495.600 94.160 ;
        RECT 4.000 91.480 496.000 92.800 ;
        RECT 4.000 90.800 495.600 91.480 ;
        RECT 4.400 90.080 495.600 90.800 ;
        RECT 4.400 89.400 496.000 90.080 ;
        RECT 4.000 88.760 496.000 89.400 ;
        RECT 4.000 87.360 495.600 88.760 ;
        RECT 4.000 86.040 496.000 87.360 ;
        RECT 4.400 84.640 495.600 86.040 ;
        RECT 4.000 83.320 496.000 84.640 ;
        RECT 4.000 81.920 495.600 83.320 ;
        RECT 4.000 81.280 496.000 81.920 ;
        RECT 4.400 80.600 496.000 81.280 ;
        RECT 4.400 79.880 495.600 80.600 ;
        RECT 4.000 79.200 495.600 79.880 ;
        RECT 4.000 77.880 496.000 79.200 ;
        RECT 4.000 76.520 495.600 77.880 ;
        RECT 4.400 76.480 495.600 76.520 ;
        RECT 4.400 75.160 496.000 76.480 ;
        RECT 4.400 75.120 495.600 75.160 ;
        RECT 4.000 73.760 495.600 75.120 ;
        RECT 4.000 72.440 496.000 73.760 ;
        RECT 4.000 71.760 495.600 72.440 ;
        RECT 4.400 71.040 495.600 71.760 ;
        RECT 4.400 70.360 496.000 71.040 ;
        RECT 4.000 69.720 496.000 70.360 ;
        RECT 4.000 68.320 495.600 69.720 ;
        RECT 4.000 67.000 496.000 68.320 ;
        RECT 4.400 65.600 495.600 67.000 ;
        RECT 4.000 64.280 496.000 65.600 ;
        RECT 4.000 62.880 495.600 64.280 ;
        RECT 4.000 62.240 496.000 62.880 ;
        RECT 4.400 61.560 496.000 62.240 ;
        RECT 4.400 60.840 495.600 61.560 ;
        RECT 4.000 60.160 495.600 60.840 ;
        RECT 4.000 58.840 496.000 60.160 ;
        RECT 4.000 57.480 495.600 58.840 ;
        RECT 4.400 57.440 495.600 57.480 ;
        RECT 4.400 56.120 496.000 57.440 ;
        RECT 4.400 56.080 495.600 56.120 ;
        RECT 4.000 54.720 495.600 56.080 ;
        RECT 4.000 53.400 496.000 54.720 ;
        RECT 4.000 52.720 495.600 53.400 ;
        RECT 4.400 52.000 495.600 52.720 ;
        RECT 4.400 51.320 496.000 52.000 ;
        RECT 4.000 50.680 496.000 51.320 ;
        RECT 4.000 49.280 495.600 50.680 ;
        RECT 4.000 47.960 496.000 49.280 ;
        RECT 4.400 46.560 495.600 47.960 ;
        RECT 4.000 45.240 496.000 46.560 ;
        RECT 4.000 43.840 495.600 45.240 ;
        RECT 4.000 43.200 496.000 43.840 ;
        RECT 4.400 42.520 496.000 43.200 ;
        RECT 4.400 41.800 495.600 42.520 ;
        RECT 4.000 41.120 495.600 41.800 ;
        RECT 4.000 39.800 496.000 41.120 ;
        RECT 4.000 38.440 495.600 39.800 ;
        RECT 4.400 38.400 495.600 38.440 ;
        RECT 4.400 37.080 496.000 38.400 ;
        RECT 4.400 37.040 495.600 37.080 ;
        RECT 4.000 35.680 495.600 37.040 ;
        RECT 4.000 33.680 496.000 35.680 ;
        RECT 4.400 32.280 496.000 33.680 ;
        RECT 4.000 28.920 496.000 32.280 ;
        RECT 4.400 27.520 496.000 28.920 ;
        RECT 4.000 24.160 496.000 27.520 ;
        RECT 4.400 22.760 496.000 24.160 ;
        RECT 4.000 19.400 496.000 22.760 ;
        RECT 4.400 18.000 496.000 19.400 ;
        RECT 4.000 14.640 496.000 18.000 ;
        RECT 4.400 13.240 496.000 14.640 ;
        RECT 4.000 6.295 496.000 13.240 ;
      LAYER met4 ;
        RECT 9.495 10.240 20.640 313.985 ;
        RECT 23.040 10.240 97.440 313.985 ;
        RECT 99.840 10.240 174.240 313.985 ;
        RECT 176.640 10.240 251.040 313.985 ;
        RECT 253.440 10.240 327.840 313.985 ;
        RECT 330.240 10.240 404.640 313.985 ;
        RECT 407.040 10.240 438.545 313.985 ;
        RECT 9.495 6.295 438.545 10.240 ;
  END
END cawb
END LIBRARY

