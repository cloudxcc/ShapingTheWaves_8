magic
tech sky130A
magscale 1 2
timestamp 1670655912
<< obsli1 >>
rect 68704 22159 528448 692753
<< obsm1 >>
rect 566 8 583450 700664
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583444 703610
rect 572 536 583444 703464
rect 710 2 1590 536
rect 1814 2 2786 536
rect 3010 2 3982 536
rect 4206 2 5178 536
rect 5402 2 6374 536
rect 6598 2 7570 536
rect 7794 2 8674 536
rect 8898 2 9870 536
rect 10094 2 11066 536
rect 11290 2 12262 536
rect 12486 2 13458 536
rect 13682 2 14654 536
rect 14878 2 15850 536
rect 16074 2 16954 536
rect 17178 2 18150 536
rect 18374 2 19346 536
rect 19570 2 20542 536
rect 20766 2 21738 536
rect 21962 2 22934 536
rect 23158 2 24130 536
rect 24354 2 25234 536
rect 25458 2 26430 536
rect 26654 2 27626 536
rect 27850 2 28822 536
rect 29046 2 30018 536
rect 30242 2 31214 536
rect 31438 2 32318 536
rect 32542 2 33514 536
rect 33738 2 34710 536
rect 34934 2 35906 536
rect 36130 2 37102 536
rect 37326 2 38298 536
rect 38522 2 39494 536
rect 39718 2 40598 536
rect 40822 2 41794 536
rect 42018 2 42990 536
rect 43214 2 44186 536
rect 44410 2 45382 536
rect 45606 2 46578 536
rect 46802 2 47774 536
rect 47998 2 48878 536
rect 49102 2 50074 536
rect 50298 2 51270 536
rect 51494 2 52466 536
rect 52690 2 53662 536
rect 53886 2 54858 536
rect 55082 2 55962 536
rect 56186 2 57158 536
rect 57382 2 58354 536
rect 58578 2 59550 536
rect 59774 2 60746 536
rect 60970 2 61942 536
rect 62166 2 63138 536
rect 63362 2 64242 536
rect 64466 2 65438 536
rect 65662 2 66634 536
rect 66858 2 67830 536
rect 68054 2 69026 536
rect 69250 2 70222 536
rect 70446 2 71418 536
rect 71642 2 72522 536
rect 72746 2 73718 536
rect 73942 2 74914 536
rect 75138 2 76110 536
rect 76334 2 77306 536
rect 77530 2 78502 536
rect 78726 2 79606 536
rect 79830 2 80802 536
rect 81026 2 81998 536
rect 82222 2 83194 536
rect 83418 2 84390 536
rect 84614 2 85586 536
rect 85810 2 86782 536
rect 87006 2 87886 536
rect 88110 2 89082 536
rect 89306 2 90278 536
rect 90502 2 91474 536
rect 91698 2 92670 536
rect 92894 2 93866 536
rect 94090 2 95062 536
rect 95286 2 96166 536
rect 96390 2 97362 536
rect 97586 2 98558 536
rect 98782 2 99754 536
rect 99978 2 100950 536
rect 101174 2 102146 536
rect 102370 2 103250 536
rect 103474 2 104446 536
rect 104670 2 105642 536
rect 105866 2 106838 536
rect 107062 2 108034 536
rect 108258 2 109230 536
rect 109454 2 110426 536
rect 110650 2 111530 536
rect 111754 2 112726 536
rect 112950 2 113922 536
rect 114146 2 115118 536
rect 115342 2 116314 536
rect 116538 2 117510 536
rect 117734 2 118706 536
rect 118930 2 119810 536
rect 120034 2 121006 536
rect 121230 2 122202 536
rect 122426 2 123398 536
rect 123622 2 124594 536
rect 124818 2 125790 536
rect 126014 2 126894 536
rect 127118 2 128090 536
rect 128314 2 129286 536
rect 129510 2 130482 536
rect 130706 2 131678 536
rect 131902 2 132874 536
rect 133098 2 134070 536
rect 134294 2 135174 536
rect 135398 2 136370 536
rect 136594 2 137566 536
rect 137790 2 138762 536
rect 138986 2 139958 536
rect 140182 2 141154 536
rect 141378 2 142350 536
rect 142574 2 143454 536
rect 143678 2 144650 536
rect 144874 2 145846 536
rect 146070 2 147042 536
rect 147266 2 148238 536
rect 148462 2 149434 536
rect 149658 2 150538 536
rect 150762 2 151734 536
rect 151958 2 152930 536
rect 153154 2 154126 536
rect 154350 2 155322 536
rect 155546 2 156518 536
rect 156742 2 157714 536
rect 157938 2 158818 536
rect 159042 2 160014 536
rect 160238 2 161210 536
rect 161434 2 162406 536
rect 162630 2 163602 536
rect 163826 2 164798 536
rect 165022 2 165994 536
rect 166218 2 167098 536
rect 167322 2 168294 536
rect 168518 2 169490 536
rect 169714 2 170686 536
rect 170910 2 171882 536
rect 172106 2 173078 536
rect 173302 2 174182 536
rect 174406 2 175378 536
rect 175602 2 176574 536
rect 176798 2 177770 536
rect 177994 2 178966 536
rect 179190 2 180162 536
rect 180386 2 181358 536
rect 181582 2 182462 536
rect 182686 2 183658 536
rect 183882 2 184854 536
rect 185078 2 186050 536
rect 186274 2 187246 536
rect 187470 2 188442 536
rect 188666 2 189638 536
rect 189862 2 190742 536
rect 190966 2 191938 536
rect 192162 2 193134 536
rect 193358 2 194330 536
rect 194554 2 195526 536
rect 195750 2 196722 536
rect 196946 2 197826 536
rect 198050 2 199022 536
rect 199246 2 200218 536
rect 200442 2 201414 536
rect 201638 2 202610 536
rect 202834 2 203806 536
rect 204030 2 205002 536
rect 205226 2 206106 536
rect 206330 2 207302 536
rect 207526 2 208498 536
rect 208722 2 209694 536
rect 209918 2 210890 536
rect 211114 2 212086 536
rect 212310 2 213282 536
rect 213506 2 214386 536
rect 214610 2 215582 536
rect 215806 2 216778 536
rect 217002 2 217974 536
rect 218198 2 219170 536
rect 219394 2 220366 536
rect 220590 2 221470 536
rect 221694 2 222666 536
rect 222890 2 223862 536
rect 224086 2 225058 536
rect 225282 2 226254 536
rect 226478 2 227450 536
rect 227674 2 228646 536
rect 228870 2 229750 536
rect 229974 2 230946 536
rect 231170 2 232142 536
rect 232366 2 233338 536
rect 233562 2 234534 536
rect 234758 2 235730 536
rect 235954 2 236926 536
rect 237150 2 238030 536
rect 238254 2 239226 536
rect 239450 2 240422 536
rect 240646 2 241618 536
rect 241842 2 242814 536
rect 243038 2 244010 536
rect 244234 2 245114 536
rect 245338 2 246310 536
rect 246534 2 247506 536
rect 247730 2 248702 536
rect 248926 2 249898 536
rect 250122 2 251094 536
rect 251318 2 252290 536
rect 252514 2 253394 536
rect 253618 2 254590 536
rect 254814 2 255786 536
rect 256010 2 256982 536
rect 257206 2 258178 536
rect 258402 2 259374 536
rect 259598 2 260570 536
rect 260794 2 261674 536
rect 261898 2 262870 536
rect 263094 2 264066 536
rect 264290 2 265262 536
rect 265486 2 266458 536
rect 266682 2 267654 536
rect 267878 2 268758 536
rect 268982 2 269954 536
rect 270178 2 271150 536
rect 271374 2 272346 536
rect 272570 2 273542 536
rect 273766 2 274738 536
rect 274962 2 275934 536
rect 276158 2 277038 536
rect 277262 2 278234 536
rect 278458 2 279430 536
rect 279654 2 280626 536
rect 280850 2 281822 536
rect 282046 2 283018 536
rect 283242 2 284214 536
rect 284438 2 285318 536
rect 285542 2 286514 536
rect 286738 2 287710 536
rect 287934 2 288906 536
rect 289130 2 290102 536
rect 290326 2 291298 536
rect 291522 2 292494 536
rect 292718 2 293598 536
rect 293822 2 294794 536
rect 295018 2 295990 536
rect 296214 2 297186 536
rect 297410 2 298382 536
rect 298606 2 299578 536
rect 299802 2 300682 536
rect 300906 2 301878 536
rect 302102 2 303074 536
rect 303298 2 304270 536
rect 304494 2 305466 536
rect 305690 2 306662 536
rect 306886 2 307858 536
rect 308082 2 308962 536
rect 309186 2 310158 536
rect 310382 2 311354 536
rect 311578 2 312550 536
rect 312774 2 313746 536
rect 313970 2 314942 536
rect 315166 2 316138 536
rect 316362 2 317242 536
rect 317466 2 318438 536
rect 318662 2 319634 536
rect 319858 2 320830 536
rect 321054 2 322026 536
rect 322250 2 323222 536
rect 323446 2 324326 536
rect 324550 2 325522 536
rect 325746 2 326718 536
rect 326942 2 327914 536
rect 328138 2 329110 536
rect 329334 2 330306 536
rect 330530 2 331502 536
rect 331726 2 332606 536
rect 332830 2 333802 536
rect 334026 2 334998 536
rect 335222 2 336194 536
rect 336418 2 337390 536
rect 337614 2 338586 536
rect 338810 2 339782 536
rect 340006 2 340886 536
rect 341110 2 342082 536
rect 342306 2 343278 536
rect 343502 2 344474 536
rect 344698 2 345670 536
rect 345894 2 346866 536
rect 347090 2 347970 536
rect 348194 2 349166 536
rect 349390 2 350362 536
rect 350586 2 351558 536
rect 351782 2 352754 536
rect 352978 2 353950 536
rect 354174 2 355146 536
rect 355370 2 356250 536
rect 356474 2 357446 536
rect 357670 2 358642 536
rect 358866 2 359838 536
rect 360062 2 361034 536
rect 361258 2 362230 536
rect 362454 2 363426 536
rect 363650 2 364530 536
rect 364754 2 365726 536
rect 365950 2 366922 536
rect 367146 2 368118 536
rect 368342 2 369314 536
rect 369538 2 370510 536
rect 370734 2 371614 536
rect 371838 2 372810 536
rect 373034 2 374006 536
rect 374230 2 375202 536
rect 375426 2 376398 536
rect 376622 2 377594 536
rect 377818 2 378790 536
rect 379014 2 379894 536
rect 380118 2 381090 536
rect 381314 2 382286 536
rect 382510 2 383482 536
rect 383706 2 384678 536
rect 384902 2 385874 536
rect 386098 2 387070 536
rect 387294 2 388174 536
rect 388398 2 389370 536
rect 389594 2 390566 536
rect 390790 2 391762 536
rect 391986 2 392958 536
rect 393182 2 394154 536
rect 394378 2 395258 536
rect 395482 2 396454 536
rect 396678 2 397650 536
rect 397874 2 398846 536
rect 399070 2 400042 536
rect 400266 2 401238 536
rect 401462 2 402434 536
rect 402658 2 403538 536
rect 403762 2 404734 536
rect 404958 2 405930 536
rect 406154 2 407126 536
rect 407350 2 408322 536
rect 408546 2 409518 536
rect 409742 2 410714 536
rect 410938 2 411818 536
rect 412042 2 413014 536
rect 413238 2 414210 536
rect 414434 2 415406 536
rect 415630 2 416602 536
rect 416826 2 417798 536
rect 418022 2 418902 536
rect 419126 2 420098 536
rect 420322 2 421294 536
rect 421518 2 422490 536
rect 422714 2 423686 536
rect 423910 2 424882 536
rect 425106 2 426078 536
rect 426302 2 427182 536
rect 427406 2 428378 536
rect 428602 2 429574 536
rect 429798 2 430770 536
rect 430994 2 431966 536
rect 432190 2 433162 536
rect 433386 2 434358 536
rect 434582 2 435462 536
rect 435686 2 436658 536
rect 436882 2 437854 536
rect 438078 2 439050 536
rect 439274 2 440246 536
rect 440470 2 441442 536
rect 441666 2 442546 536
rect 442770 2 443742 536
rect 443966 2 444938 536
rect 445162 2 446134 536
rect 446358 2 447330 536
rect 447554 2 448526 536
rect 448750 2 449722 536
rect 449946 2 450826 536
rect 451050 2 452022 536
rect 452246 2 453218 536
rect 453442 2 454414 536
rect 454638 2 455610 536
rect 455834 2 456806 536
rect 457030 2 458002 536
rect 458226 2 459106 536
rect 459330 2 460302 536
rect 460526 2 461498 536
rect 461722 2 462694 536
rect 462918 2 463890 536
rect 464114 2 465086 536
rect 465310 2 466190 536
rect 466414 2 467386 536
rect 467610 2 468582 536
rect 468806 2 469778 536
rect 470002 2 470974 536
rect 471198 2 472170 536
rect 472394 2 473366 536
rect 473590 2 474470 536
rect 474694 2 475666 536
rect 475890 2 476862 536
rect 477086 2 478058 536
rect 478282 2 479254 536
rect 479478 2 480450 536
rect 480674 2 481646 536
rect 481870 2 482750 536
rect 482974 2 483946 536
rect 484170 2 485142 536
rect 485366 2 486338 536
rect 486562 2 487534 536
rect 487758 2 488730 536
rect 488954 2 489834 536
rect 490058 2 491030 536
rect 491254 2 492226 536
rect 492450 2 493422 536
rect 493646 2 494618 536
rect 494842 2 495814 536
rect 496038 2 497010 536
rect 497234 2 498114 536
rect 498338 2 499310 536
rect 499534 2 500506 536
rect 500730 2 501702 536
rect 501926 2 502898 536
rect 503122 2 504094 536
rect 504318 2 505290 536
rect 505514 2 506394 536
rect 506618 2 507590 536
rect 507814 2 508786 536
rect 509010 2 509982 536
rect 510206 2 511178 536
rect 511402 2 512374 536
rect 512598 2 513478 536
rect 513702 2 514674 536
rect 514898 2 515870 536
rect 516094 2 517066 536
rect 517290 2 518262 536
rect 518486 2 519458 536
rect 519682 2 520654 536
rect 520878 2 521758 536
rect 521982 2 522954 536
rect 523178 2 524150 536
rect 524374 2 525346 536
rect 525570 2 526542 536
rect 526766 2 527738 536
rect 527962 2 528934 536
rect 529158 2 530038 536
rect 530262 2 531234 536
rect 531458 2 532430 536
rect 532654 2 533626 536
rect 533850 2 534822 536
rect 535046 2 536018 536
rect 536242 2 537122 536
rect 537346 2 538318 536
rect 538542 2 539514 536
rect 539738 2 540710 536
rect 540934 2 541906 536
rect 542130 2 543102 536
rect 543326 2 544298 536
rect 544522 2 545402 536
rect 545626 2 546598 536
rect 546822 2 547794 536
rect 548018 2 548990 536
rect 549214 2 550186 536
rect 550410 2 551382 536
rect 551606 2 552578 536
rect 552802 2 553682 536
rect 553906 2 554878 536
rect 555102 2 556074 536
rect 556298 2 557270 536
rect 557494 2 558466 536
rect 558690 2 559662 536
rect 559886 2 560766 536
rect 560990 2 561962 536
rect 562186 2 563158 536
rect 563382 2 564354 536
rect 564578 2 565550 536
rect 565774 2 566746 536
rect 566970 2 567942 536
rect 568166 2 569046 536
rect 569270 2 570242 536
rect 570466 2 571438 536
rect 571662 2 572634 536
rect 572858 2 573830 536
rect 574054 2 575026 536
rect 575250 2 576222 536
rect 576446 2 577326 536
rect 577550 2 578522 536
rect 578746 2 579718 536
rect 579942 2 580914 536
rect 581138 2 582110 536
rect 582334 2 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583520 700365
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 35 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 5514 -7654 6134 711590
rect 9234 -7654 9854 711590
rect 12954 -7654 13574 711590
rect 16674 -7654 17294 711590
rect 20394 -7654 21014 711590
rect 24114 -7654 24734 711590
rect 27834 -7654 28454 711590
rect 31794 -7654 32414 711590
rect 35514 -7654 36134 711590
rect 39234 654660 39854 711590
rect 42954 654660 43574 711590
rect 46674 654660 47294 711590
rect 50394 654660 51014 711590
rect 54114 654660 54734 711590
rect 57834 654660 58454 711590
rect 61794 654660 62414 711590
rect 65514 654660 66134 711590
rect 69234 654784 69854 711590
rect 72954 654784 73574 711590
rect 76674 654784 77294 711590
rect 80394 654784 81014 711590
rect 84114 654784 84734 711590
rect 87834 654784 88454 711590
rect 91794 654784 92414 711590
rect 95514 654784 96134 711590
rect 99234 654784 99854 711590
rect 102954 654784 103574 711590
rect 106674 654784 107294 711590
rect 110394 654660 111014 711590
rect 114114 654660 114734 711590
rect 117834 654660 118454 711590
rect 121794 654784 122414 711590
rect 125514 654660 126134 711590
rect 129234 654660 129854 711590
rect 132954 654660 133574 711590
rect 136674 654660 137294 711590
rect 39234 508660 39854 570064
rect 42954 508660 43574 570064
rect 46674 508660 47294 570064
rect 50394 508660 51014 570064
rect 54114 508660 54734 570064
rect 57834 508660 58454 569940
rect 61794 508660 62414 569940
rect 65514 508660 66134 570064
rect 69234 508784 69854 569940
rect 72954 508784 73574 569940
rect 76674 508784 77294 569940
rect 80394 508784 81014 569940
rect 84114 508784 84734 569940
rect 87834 508784 88454 569940
rect 91794 508784 92414 569940
rect 95514 508784 96134 569940
rect 99234 508784 99854 569940
rect 102954 508784 103574 569940
rect 106674 508784 107294 569940
rect 110394 508660 111014 570064
rect 114114 508660 114734 570064
rect 117834 508660 118454 570064
rect 121794 508784 122414 570064
rect 125514 508660 126134 569940
rect 129234 508660 129854 570064
rect 132954 508660 133574 570064
rect 136674 508660 137294 570064
rect 50394 378660 51014 424064
rect 54114 378660 54734 424064
rect 57834 378660 58454 423940
rect 61794 378660 62414 423940
rect 69234 378784 69854 423940
rect 72954 378784 73574 423940
rect 76674 378784 77294 423940
rect 80394 378784 81014 423940
rect 84114 378784 84734 423940
rect 87834 378784 88454 423940
rect 91794 378784 92414 423940
rect 95514 378784 96134 423940
rect 99234 378784 99854 423940
rect 102954 378784 103574 423940
rect 106674 378784 107294 423940
rect 110394 378660 111014 424064
rect 114114 378660 114734 424064
rect 117834 378660 118454 424064
rect 121794 378784 122414 424064
rect 39234 240660 39854 294064
rect 42954 240660 43574 294064
rect 46674 240660 47294 294064
rect 50394 240660 51014 294064
rect 61794 240660 62414 293940
rect 65514 240660 66134 294064
rect 69234 240784 69854 293940
rect 72954 240784 73574 293940
rect 76674 240784 77294 293940
rect 80394 240784 81014 293940
rect 84114 240784 84734 293940
rect 87834 240784 88454 293940
rect 91794 240784 92414 293940
rect 95514 240784 96134 293940
rect 99234 240784 99854 293940
rect 102954 240784 103574 293940
rect 106674 240784 107294 293940
rect 110394 240660 111014 294064
rect 121794 240784 122414 294064
rect 125514 240660 126134 293940
rect 129234 240660 129854 294064
rect 132954 240660 133574 294064
rect 136674 240660 137294 294064
rect 42954 102660 43574 156064
rect 46674 102660 47294 156064
rect 50394 102660 51014 156064
rect 54114 102660 54734 156064
rect 57834 102660 58454 155940
rect 61794 102660 62414 155940
rect 69234 102784 69854 155940
rect 72954 102784 73574 155940
rect 76674 102784 77294 155940
rect 80394 102784 81014 155940
rect 84114 102784 84734 155940
rect 87834 102784 88454 155940
rect 91794 102784 92414 155940
rect 95514 102784 96134 155940
rect 99234 102784 99854 155940
rect 102954 102784 103574 155940
rect 106674 102784 107294 155940
rect 110394 102660 111014 156064
rect 114114 102660 114734 156064
rect 117834 102660 118454 156064
rect 121794 102784 122414 156064
rect 132954 102660 133574 156064
rect 136674 102660 137294 156064
rect 39234 -7654 39854 18064
rect 42954 -7654 43574 18064
rect 46674 -7654 47294 18064
rect 61794 -7654 62414 17940
rect 65514 -7654 66134 18064
rect 69234 -7654 69854 17940
rect 72954 -7654 73574 17940
rect 76674 -7654 77294 17940
rect 91794 -7654 92414 17940
rect 95514 -7654 96134 17940
rect 99234 -7654 99854 17940
rect 102954 -7654 103574 17940
rect 106674 -7654 107294 17940
rect 121794 -7654 122414 18064
rect 125514 -7654 126134 17940
rect 129234 -7654 129854 18064
rect 132954 -7654 133574 18064
rect 136674 -7654 137294 18064
rect 140394 -7654 141014 711590
rect 144114 -7654 144734 711590
rect 147834 -7654 148454 711590
rect 151794 -7654 152414 711590
rect 155514 -7654 156134 711590
rect 159234 -7654 159854 711590
rect 162954 -7654 163574 711590
rect 166674 -7654 167294 711590
rect 170394 -7654 171014 711590
rect 174114 -7654 174734 711590
rect 177834 654660 178454 711590
rect 181794 654660 182414 711590
rect 185514 654660 186134 711590
rect 189234 654660 189854 711590
rect 192954 654660 193574 711590
rect 196674 654660 197294 711590
rect 200394 654660 201014 711590
rect 204114 654660 204734 711590
rect 207834 654660 208454 711590
rect 215514 654784 216134 711590
rect 219234 654784 219854 711590
rect 222954 654784 223574 711590
rect 230394 654784 231014 711590
rect 234114 654784 234734 711590
rect 237834 654784 238454 711590
rect 241794 654784 242414 711590
rect 245514 654784 246134 711590
rect 249234 654660 249854 711590
rect 252954 654660 253574 711590
rect 256674 654660 257294 711590
rect 260394 654660 261014 711590
rect 264114 654660 264734 711590
rect 267834 654660 268454 711590
rect 271794 654784 272414 711590
rect 275514 654660 276134 711590
rect 279234 654660 279854 711590
rect 177834 -7654 178454 570064
rect 207834 539417 208454 570064
rect 237834 539417 238454 569940
rect 267834 539417 268454 570064
rect 282954 539417 283574 711590
rect 286674 539417 287294 711590
rect 290394 539417 291014 711590
rect 294114 539417 294734 711590
rect 297834 539417 298454 711590
rect 301794 539417 302414 711590
rect 305514 539417 306134 711590
rect 309234 539417 309854 711590
rect 312954 539417 313574 711590
rect 316674 539417 317294 711590
rect 320394 654784 321014 711590
rect 324114 654660 324734 711590
rect 327834 654660 328454 711590
rect 331794 654660 332414 711590
rect 335514 654660 336134 711590
rect 339234 654660 339854 711590
rect 342954 654660 343574 711590
rect 346674 654660 347294 711590
rect 350394 654784 351014 711590
rect 354114 654784 354734 711590
rect 357834 654784 358454 711590
rect 361794 654784 362414 711590
rect 365514 654784 366134 711590
rect 369234 654784 369854 711590
rect 372954 654784 373574 711590
rect 376674 654784 377294 711590
rect 380394 654784 381014 711590
rect 384114 654784 384734 711590
rect 387834 654784 388454 711590
rect 391794 654660 392414 711590
rect 395514 654660 396134 711590
rect 399234 654660 399854 711590
rect 402954 654660 403574 711590
rect 406674 654660 407294 711590
rect 410394 654660 411014 711590
rect 414114 654660 414734 711590
rect 417834 654784 418454 711590
rect 327834 539417 328454 570064
rect 357834 539417 358454 569940
rect 387834 539417 388454 569940
rect 417834 539417 418454 569940
rect 181794 84857 182414 140559
rect 185514 84857 186134 140559
rect 189234 84857 189854 140559
rect 192954 84857 193574 140559
rect 196674 84857 197294 140559
rect 204114 84857 204734 140559
rect 207834 84857 208454 140559
rect 211794 84857 212414 140559
rect 215514 84857 216134 140559
rect 219234 84857 219854 140559
rect 222954 84857 223574 140559
rect 226674 84857 227294 140559
rect 234114 84857 234734 140559
rect 237834 84857 238454 140559
rect 241794 84857 242414 140559
rect 249234 84857 249854 140559
rect 252954 84857 253574 140559
rect 256674 84857 257294 140559
rect 264114 84857 264734 140559
rect 267834 84857 268454 140559
rect 181794 -7654 182414 19199
rect 185514 -7654 186134 19199
rect 189234 -7654 189854 19199
rect 192954 -7654 193574 19199
rect 196674 -7654 197294 19199
rect 211794 -7654 212414 19199
rect 215514 -7654 216134 19199
rect 219234 -7654 219854 19199
rect 222954 -7654 223574 19199
rect 226674 -7654 227294 19199
rect 241794 -7654 242414 19199
rect 245514 -7654 246134 19199
rect 249234 -7654 249854 19199
rect 252954 -7654 253574 19199
rect 256674 -7654 257294 19199
rect 271794 -7654 272414 140559
rect 275514 -7654 276134 140559
rect 279234 -7654 279854 140559
rect 282954 -7654 283574 140559
rect 286674 -7654 287294 140559
rect 290394 -7654 291014 140559
rect 294114 -7654 294734 140559
rect 297834 -7654 298454 140559
rect 301794 -7654 302414 140559
rect 305514 -7654 306134 140559
rect 309234 -7654 309854 140559
rect 312954 -7654 313574 140559
rect 316674 -7654 317294 140559
rect 342954 102660 343574 140559
rect 346674 102660 347294 140559
rect 372954 102784 373574 140559
rect 376674 102784 377294 140559
rect 402954 102784 403574 140559
rect 406674 102660 407294 140559
rect 331794 -7654 332414 18064
rect 335514 -7654 336134 18064
rect 339234 -7654 339854 18064
rect 342954 -7654 343574 18064
rect 346674 -7654 347294 18064
rect 361794 -7654 362414 18064
rect 365514 -7654 366134 17940
rect 369234 -7654 369854 17940
rect 372954 -7654 373574 17940
rect 376674 -7654 377294 17940
rect 391794 -7654 392414 18064
rect 395514 -7654 396134 18064
rect 399234 -7654 399854 18064
rect 402954 -7654 403574 18064
rect 406674 -7654 407294 18064
rect 421794 -7654 422414 711590
rect 425514 -7654 426134 711590
rect 429234 -7654 429854 711590
rect 432954 -7654 433574 711590
rect 436674 -7654 437294 711590
rect 440394 -7654 441014 711590
rect 444114 -7654 444734 711590
rect 447834 -7654 448454 711590
rect 451794 -7654 452414 711590
rect 455514 -7654 456134 711590
rect 459234 654660 459854 711590
rect 462954 654660 463574 711590
rect 466674 654660 467294 711590
rect 470394 654660 471014 711590
rect 474114 654660 474734 711590
rect 477834 654660 478454 711590
rect 481794 654660 482414 711590
rect 485514 654660 486134 711590
rect 489234 654784 489854 711590
rect 492954 654784 493574 711590
rect 496674 654784 497294 711590
rect 500394 654784 501014 711590
rect 504114 654784 504734 711590
rect 507834 654784 508454 711590
rect 511794 654784 512414 711590
rect 515514 654784 516134 711590
rect 519234 654784 519854 711590
rect 522954 654784 523574 711590
rect 526674 654784 527294 711590
rect 530394 654660 531014 711590
rect 534114 654660 534734 711590
rect 537834 654660 538454 711590
rect 541794 654784 542414 711590
rect 545514 654660 546134 711590
rect 549234 654660 549854 711590
rect 552954 654660 553574 711590
rect 556674 654660 557294 711590
rect 459234 508660 459854 570064
rect 462954 508660 463574 570064
rect 466674 508660 467294 570064
rect 470394 508660 471014 570064
rect 474114 508660 474734 570064
rect 477834 508660 478454 569940
rect 481794 508660 482414 569940
rect 485514 508660 486134 570064
rect 489234 508784 489854 569940
rect 492954 508784 493574 569940
rect 496674 508784 497294 569940
rect 500394 508784 501014 569940
rect 504114 508784 504734 569940
rect 507834 508784 508454 569940
rect 511794 508784 512414 569940
rect 515514 508784 516134 569940
rect 519234 508784 519854 569940
rect 522954 508784 523574 569940
rect 526674 508784 527294 569940
rect 530394 508660 531014 570064
rect 534114 508660 534734 570064
rect 537834 508660 538454 570064
rect 541794 508784 542414 570064
rect 545514 508660 546134 569940
rect 549234 508660 549854 570064
rect 552954 508660 553574 570064
rect 556674 508660 557294 570064
rect 470394 378660 471014 424064
rect 474114 378660 474734 424064
rect 477834 378660 478454 423940
rect 481794 378660 482414 423940
rect 489234 378784 489854 423940
rect 492954 378784 493574 423940
rect 496674 378784 497294 423940
rect 500394 378784 501014 423940
rect 504114 378784 504734 423940
rect 507834 378784 508454 423940
rect 511794 378784 512414 423940
rect 515514 378784 516134 423940
rect 519234 378784 519854 423940
rect 522954 378784 523574 423940
rect 526674 378784 527294 423940
rect 530394 378660 531014 424064
rect 534114 378660 534734 424064
rect 537834 378660 538454 424064
rect 541794 378784 542414 424064
rect 459234 240660 459854 294064
rect 462954 240660 463574 294064
rect 466674 240660 467294 294064
rect 470394 240660 471014 294064
rect 481794 240660 482414 293940
rect 485514 240660 486134 294064
rect 489234 240784 489854 293940
rect 492954 240784 493574 293940
rect 496674 240784 497294 293940
rect 500394 240784 501014 293940
rect 504114 240784 504734 293940
rect 507834 240784 508454 293940
rect 511794 240784 512414 293940
rect 515514 240784 516134 293940
rect 519234 240784 519854 293940
rect 522954 240784 523574 293940
rect 526674 240784 527294 293940
rect 530394 240660 531014 294064
rect 541794 240784 542414 294064
rect 545514 240660 546134 293940
rect 549234 240660 549854 294064
rect 552954 240660 553574 294064
rect 556674 240660 557294 294064
rect 462954 102660 463574 156064
rect 466674 102660 467294 156064
rect 470394 102660 471014 156064
rect 474114 102660 474734 156064
rect 477834 102660 478454 155940
rect 481794 102660 482414 155940
rect 489234 102784 489854 155940
rect 492954 102784 493574 155940
rect 496674 102784 497294 155940
rect 500394 102784 501014 155940
rect 504114 102784 504734 155940
rect 507834 102784 508454 155940
rect 511794 102784 512414 155940
rect 515514 102784 516134 155940
rect 519234 102784 519854 155940
rect 522954 102784 523574 155940
rect 526674 102784 527294 155940
rect 530394 102660 531014 156064
rect 534114 102660 534734 156064
rect 537834 102660 538454 156064
rect 541794 102784 542414 156064
rect 552954 102660 553574 156064
rect 556674 102660 557294 156064
rect 459234 -7654 459854 18064
rect 462954 -7654 463574 18064
rect 466674 -7654 467294 18064
rect 481794 -7654 482414 17940
rect 485514 -7654 486134 18064
rect 489234 -7654 489854 17940
rect 492954 -7654 493574 17940
rect 496674 -7654 497294 17940
rect 511794 -7654 512414 17940
rect 515514 -7654 516134 17940
rect 519234 -7654 519854 17940
rect 522954 -7654 523574 17940
rect 526674 -7654 527294 17940
rect 541794 -7654 542414 18064
rect 545514 -7654 546134 17940
rect 549234 -7654 549854 18064
rect 552954 -7654 553574 18064
rect 556674 -7654 557294 18064
rect 560394 -7654 561014 711590
rect 564114 -7654 564734 711590
rect 567834 -7654 568454 711590
rect 571794 -7654 572414 711590
rect 575514 -7654 576134 711590
rect 579234 -7654 579854 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 40000 654580 42874 700365
rect 43654 654580 46594 700365
rect 47374 654580 50314 700365
rect 51094 654580 54034 700365
rect 54814 654580 57754 700365
rect 58534 654580 61714 700365
rect 62494 654580 65434 700365
rect 66214 654704 69154 700365
rect 69934 654704 72874 700365
rect 73654 654704 76594 700365
rect 77374 654704 80314 700365
rect 81094 654704 84034 700365
rect 84814 654704 87754 700365
rect 88534 654704 91714 700365
rect 92494 654704 95434 700365
rect 96214 654704 99154 700365
rect 99934 654704 102874 700365
rect 103654 654704 106594 700365
rect 107374 654704 110314 700365
rect 66214 654580 110314 654704
rect 111094 654580 114034 700365
rect 114814 654580 117754 700365
rect 118534 654704 121714 700365
rect 122494 654704 125434 700365
rect 118534 654580 125434 654704
rect 126214 654580 129154 700365
rect 129934 654580 132874 700365
rect 133654 654580 136594 700365
rect 137374 654580 140314 700365
rect 40000 570144 140314 654580
rect 40000 508580 42874 570144
rect 43654 508580 46594 570144
rect 47374 508580 50314 570144
rect 51094 508580 54034 570144
rect 54814 570020 65434 570144
rect 54814 508580 57754 570020
rect 58534 508580 61714 570020
rect 62494 508580 65434 570020
rect 66214 570020 110314 570144
rect 66214 508704 69154 570020
rect 69934 508704 72874 570020
rect 73654 508704 76594 570020
rect 77374 508704 80314 570020
rect 81094 508704 84034 570020
rect 84814 508704 87754 570020
rect 88534 508704 91714 570020
rect 92494 508704 95434 570020
rect 96214 508704 99154 570020
rect 99934 508704 102874 570020
rect 103654 508704 106594 570020
rect 107374 508704 110314 570020
rect 66214 508580 110314 508704
rect 111094 508580 114034 570144
rect 114814 508580 117754 570144
rect 118534 508704 121714 570144
rect 122494 570020 129154 570144
rect 122494 508704 125434 570020
rect 118534 508580 125434 508704
rect 126214 508580 129154 570020
rect 129934 508580 132874 570144
rect 133654 508580 136594 570144
rect 137374 508580 140314 570144
rect 40000 424144 140314 508580
rect 40000 378580 50314 424144
rect 51094 378580 54034 424144
rect 54814 424020 110314 424144
rect 54814 378580 57754 424020
rect 58534 378580 61714 424020
rect 62494 378704 69154 424020
rect 69934 378704 72874 424020
rect 73654 378704 76594 424020
rect 77374 378704 80314 424020
rect 81094 378704 84034 424020
rect 84814 378704 87754 424020
rect 88534 378704 91714 424020
rect 92494 378704 95434 424020
rect 96214 378704 99154 424020
rect 99934 378704 102874 424020
rect 103654 378704 106594 424020
rect 107374 378704 110314 424020
rect 62494 378580 110314 378704
rect 111094 378580 114034 424144
rect 114814 378580 117754 424144
rect 118534 378704 121714 424144
rect 122494 378704 140314 424144
rect 118534 378580 140314 378704
rect 40000 294144 140314 378580
rect 40000 240580 42874 294144
rect 43654 240580 46594 294144
rect 47374 240580 50314 294144
rect 51094 294020 65434 294144
rect 51094 240580 61714 294020
rect 62494 240580 65434 294020
rect 66214 294020 110314 294144
rect 66214 240704 69154 294020
rect 69934 240704 72874 294020
rect 73654 240704 76594 294020
rect 77374 240704 80314 294020
rect 81094 240704 84034 294020
rect 84814 240704 87754 294020
rect 88534 240704 91714 294020
rect 92494 240704 95434 294020
rect 96214 240704 99154 294020
rect 99934 240704 102874 294020
rect 103654 240704 106594 294020
rect 107374 240704 110314 294020
rect 66214 240580 110314 240704
rect 111094 240704 121714 294144
rect 122494 294020 129154 294144
rect 122494 240704 125434 294020
rect 111094 240580 125434 240704
rect 126214 240580 129154 294020
rect 129934 240580 132874 294144
rect 133654 240580 136594 294144
rect 137374 240580 140314 294144
rect 40000 156144 140314 240580
rect 40000 102580 42874 156144
rect 43654 102580 46594 156144
rect 47374 102580 50314 156144
rect 51094 102580 54034 156144
rect 54814 156020 110314 156144
rect 54814 102580 57754 156020
rect 58534 102580 61714 156020
rect 62494 102704 69154 156020
rect 69934 102704 72874 156020
rect 73654 102704 76594 156020
rect 77374 102704 80314 156020
rect 81094 102704 84034 156020
rect 84814 102704 87754 156020
rect 88534 102704 91714 156020
rect 92494 102704 95434 156020
rect 96214 102704 99154 156020
rect 99934 102704 102874 156020
rect 103654 102704 106594 156020
rect 107374 102704 110314 156020
rect 62494 102580 110314 102704
rect 111094 102580 114034 156144
rect 114814 102580 117754 156144
rect 118534 102704 121714 156144
rect 122494 102704 132874 156144
rect 118534 102580 132874 102704
rect 133654 102580 136594 156144
rect 137374 102580 140314 156144
rect 40000 18144 140314 102580
rect 40000 8195 42874 18144
rect 43654 8195 46594 18144
rect 47374 18020 65434 18144
rect 47374 8195 61714 18020
rect 62494 8195 65434 18020
rect 66214 18020 121714 18144
rect 66214 8195 69154 18020
rect 69934 8195 72874 18020
rect 73654 8195 76594 18020
rect 77374 8195 91714 18020
rect 92494 8195 95434 18020
rect 96214 8195 99154 18020
rect 99934 8195 102874 18020
rect 103654 8195 106594 18020
rect 107374 8195 121714 18020
rect 122494 18020 129154 18144
rect 122494 8195 125434 18020
rect 126214 8195 129154 18020
rect 129934 8195 132874 18144
rect 133654 8195 136594 18144
rect 137374 8195 140314 18144
rect 141094 8195 144034 700365
rect 144814 8195 147754 700365
rect 148534 8195 151714 700365
rect 152494 8195 155434 700365
rect 156214 8195 159154 700365
rect 159934 8195 162874 700365
rect 163654 8195 166594 700365
rect 167374 8195 170314 700365
rect 171094 8195 174034 700365
rect 174814 654580 177754 700365
rect 178534 654580 181714 700365
rect 182494 654580 185434 700365
rect 186214 654580 189154 700365
rect 189934 654580 192874 700365
rect 193654 654580 196594 700365
rect 197374 654580 200314 700365
rect 201094 654580 204034 700365
rect 204814 654580 207754 700365
rect 208534 654704 215434 700365
rect 216214 654704 219154 700365
rect 219934 654704 222874 700365
rect 223654 654704 230314 700365
rect 231094 654704 234034 700365
rect 234814 654704 237754 700365
rect 238534 654704 241714 700365
rect 242494 654704 245434 700365
rect 246214 654704 249154 700365
rect 208534 654580 249154 654704
rect 249934 654580 252874 700365
rect 253654 654580 256594 700365
rect 257374 654580 260314 700365
rect 261094 654580 264034 700365
rect 264814 654580 267754 700365
rect 268534 654704 271714 700365
rect 272494 654704 275434 700365
rect 268534 654580 275434 654704
rect 276214 654580 279154 700365
rect 279934 654580 282874 700365
rect 174814 570144 282874 654580
rect 174814 8195 177754 570144
rect 178534 539337 207754 570144
rect 208534 570020 267754 570144
rect 208534 539337 237754 570020
rect 238534 539337 267754 570020
rect 268534 539337 282874 570144
rect 283654 539337 286594 700365
rect 287374 539337 290314 700365
rect 291094 539337 294034 700365
rect 294814 539337 297754 700365
rect 298534 539337 301714 700365
rect 302494 539337 305434 700365
rect 306214 539337 309154 700365
rect 309934 539337 312874 700365
rect 313654 539337 316594 700365
rect 317374 654704 320314 700365
rect 321094 654704 324034 700365
rect 317374 654580 324034 654704
rect 324814 654580 327754 700365
rect 328534 654580 331714 700365
rect 332494 654580 335434 700365
rect 336214 654580 339154 700365
rect 339934 654580 342874 700365
rect 343654 654580 346594 700365
rect 347374 654704 350314 700365
rect 351094 654704 354034 700365
rect 354814 654704 357754 700365
rect 358534 654704 361714 700365
rect 362494 654704 365434 700365
rect 366214 654704 369154 700365
rect 369934 654704 372874 700365
rect 373654 654704 376594 700365
rect 377374 654704 380314 700365
rect 381094 654704 384034 700365
rect 384814 654704 387754 700365
rect 388534 654704 391714 700365
rect 347374 654580 391714 654704
rect 392494 654580 395434 700365
rect 396214 654580 399154 700365
rect 399934 654580 402874 700365
rect 403654 654580 406594 700365
rect 407374 654580 410314 700365
rect 411094 654580 414034 700365
rect 414814 654704 417754 700365
rect 418534 654704 421714 700365
rect 414814 654580 421714 654704
rect 317374 570144 421714 654580
rect 317374 539337 327754 570144
rect 328534 570020 421714 570144
rect 328534 539337 357754 570020
rect 358534 539337 387754 570020
rect 388534 539337 417754 570020
rect 418534 539337 421714 570020
rect 178534 140639 421714 539337
rect 178534 84777 181714 140639
rect 182494 84777 185434 140639
rect 186214 84777 189154 140639
rect 189934 84777 192874 140639
rect 193654 84777 196594 140639
rect 197374 84777 204034 140639
rect 204814 84777 207754 140639
rect 208534 84777 211714 140639
rect 212494 84777 215434 140639
rect 216214 84777 219154 140639
rect 219934 84777 222874 140639
rect 223654 84777 226594 140639
rect 227374 84777 234034 140639
rect 234814 84777 237754 140639
rect 238534 84777 241714 140639
rect 242494 84777 249154 140639
rect 249934 84777 252874 140639
rect 253654 84777 256594 140639
rect 257374 84777 264034 140639
rect 264814 84777 267754 140639
rect 268534 84777 271714 140639
rect 178534 19279 271714 84777
rect 178534 8195 181714 19279
rect 182494 8195 185434 19279
rect 186214 8195 189154 19279
rect 189934 8195 192874 19279
rect 193654 8195 196594 19279
rect 197374 8195 211714 19279
rect 212494 8195 215434 19279
rect 216214 8195 219154 19279
rect 219934 8195 222874 19279
rect 223654 8195 226594 19279
rect 227374 8195 241714 19279
rect 242494 8195 245434 19279
rect 246214 8195 249154 19279
rect 249934 8195 252874 19279
rect 253654 8195 256594 19279
rect 257374 8195 271714 19279
rect 272494 8195 275434 140639
rect 276214 8195 279154 140639
rect 279934 8195 282874 140639
rect 283654 8195 286594 140639
rect 287374 8195 290314 140639
rect 291094 8195 294034 140639
rect 294814 8195 297754 140639
rect 298534 8195 301714 140639
rect 302494 8195 305434 140639
rect 306214 8195 309154 140639
rect 309934 8195 312874 140639
rect 313654 8195 316594 140639
rect 317374 102580 342874 140639
rect 343654 102580 346594 140639
rect 347374 102704 372874 140639
rect 373654 102704 376594 140639
rect 377374 102704 402874 140639
rect 403654 102704 406594 140639
rect 347374 102580 406594 102704
rect 407374 102580 421714 140639
rect 317374 18144 421714 102580
rect 317374 8195 331714 18144
rect 332494 8195 335434 18144
rect 336214 8195 339154 18144
rect 339934 8195 342874 18144
rect 343654 8195 346594 18144
rect 347374 8195 361714 18144
rect 362494 18020 391714 18144
rect 362494 8195 365434 18020
rect 366214 8195 369154 18020
rect 369934 8195 372874 18020
rect 373654 8195 376594 18020
rect 377374 8195 391714 18020
rect 392494 8195 395434 18144
rect 396214 8195 399154 18144
rect 399934 8195 402874 18144
rect 403654 8195 406594 18144
rect 407374 8195 421714 18144
rect 422494 8195 425434 700365
rect 426214 8195 429154 700365
rect 429934 8195 432874 700365
rect 433654 8195 436594 700365
rect 437374 8195 440314 700365
rect 441094 8195 444034 700365
rect 444814 8195 447754 700365
rect 448534 8195 451714 700365
rect 452494 8195 455434 700365
rect 456214 654580 459154 700365
rect 459934 654580 462874 700365
rect 463654 654580 466594 700365
rect 467374 654580 470314 700365
rect 471094 654580 474034 700365
rect 474814 654580 477754 700365
rect 478534 654580 481714 700365
rect 482494 654580 485434 700365
rect 486214 654704 489154 700365
rect 489934 654704 492874 700365
rect 493654 654704 496594 700365
rect 497374 654704 500314 700365
rect 501094 654704 504034 700365
rect 504814 654704 507754 700365
rect 508534 654704 511714 700365
rect 512494 654704 515434 700365
rect 516214 654704 519154 700365
rect 519934 654704 522874 700365
rect 523654 654704 526594 700365
rect 527374 654704 530314 700365
rect 486214 654580 530314 654704
rect 531094 654580 534034 700365
rect 534814 654580 537754 700365
rect 538534 654704 541714 700365
rect 542494 654704 545434 700365
rect 538534 654580 545434 654704
rect 546214 654580 549154 700365
rect 549934 654580 552874 700365
rect 553654 654580 556594 700365
rect 557374 654580 558676 700365
rect 456214 570144 558676 654580
rect 456214 508580 459154 570144
rect 459934 508580 462874 570144
rect 463654 508580 466594 570144
rect 467374 508580 470314 570144
rect 471094 508580 474034 570144
rect 474814 570020 485434 570144
rect 474814 508580 477754 570020
rect 478534 508580 481714 570020
rect 482494 508580 485434 570020
rect 486214 570020 530314 570144
rect 486214 508704 489154 570020
rect 489934 508704 492874 570020
rect 493654 508704 496594 570020
rect 497374 508704 500314 570020
rect 501094 508704 504034 570020
rect 504814 508704 507754 570020
rect 508534 508704 511714 570020
rect 512494 508704 515434 570020
rect 516214 508704 519154 570020
rect 519934 508704 522874 570020
rect 523654 508704 526594 570020
rect 527374 508704 530314 570020
rect 486214 508580 530314 508704
rect 531094 508580 534034 570144
rect 534814 508580 537754 570144
rect 538534 508704 541714 570144
rect 542494 570020 549154 570144
rect 542494 508704 545434 570020
rect 538534 508580 545434 508704
rect 546214 508580 549154 570020
rect 549934 508580 552874 570144
rect 553654 508580 556594 570144
rect 557374 508580 558676 570144
rect 456214 424144 558676 508580
rect 456214 378580 470314 424144
rect 471094 378580 474034 424144
rect 474814 424020 530314 424144
rect 474814 378580 477754 424020
rect 478534 378580 481714 424020
rect 482494 378704 489154 424020
rect 489934 378704 492874 424020
rect 493654 378704 496594 424020
rect 497374 378704 500314 424020
rect 501094 378704 504034 424020
rect 504814 378704 507754 424020
rect 508534 378704 511714 424020
rect 512494 378704 515434 424020
rect 516214 378704 519154 424020
rect 519934 378704 522874 424020
rect 523654 378704 526594 424020
rect 527374 378704 530314 424020
rect 482494 378580 530314 378704
rect 531094 378580 534034 424144
rect 534814 378580 537754 424144
rect 538534 378704 541714 424144
rect 542494 378704 558676 424144
rect 538534 378580 558676 378704
rect 456214 294144 558676 378580
rect 456214 240580 459154 294144
rect 459934 240580 462874 294144
rect 463654 240580 466594 294144
rect 467374 240580 470314 294144
rect 471094 294020 485434 294144
rect 471094 240580 481714 294020
rect 482494 240580 485434 294020
rect 486214 294020 530314 294144
rect 486214 240704 489154 294020
rect 489934 240704 492874 294020
rect 493654 240704 496594 294020
rect 497374 240704 500314 294020
rect 501094 240704 504034 294020
rect 504814 240704 507754 294020
rect 508534 240704 511714 294020
rect 512494 240704 515434 294020
rect 516214 240704 519154 294020
rect 519934 240704 522874 294020
rect 523654 240704 526594 294020
rect 527374 240704 530314 294020
rect 486214 240580 530314 240704
rect 531094 240704 541714 294144
rect 542494 294020 549154 294144
rect 542494 240704 545434 294020
rect 531094 240580 545434 240704
rect 546214 240580 549154 294020
rect 549934 240580 552874 294144
rect 553654 240580 556594 294144
rect 557374 240580 558676 294144
rect 456214 156144 558676 240580
rect 456214 102580 462874 156144
rect 463654 102580 466594 156144
rect 467374 102580 470314 156144
rect 471094 102580 474034 156144
rect 474814 156020 530314 156144
rect 474814 102580 477754 156020
rect 478534 102580 481714 156020
rect 482494 102704 489154 156020
rect 489934 102704 492874 156020
rect 493654 102704 496594 156020
rect 497374 102704 500314 156020
rect 501094 102704 504034 156020
rect 504814 102704 507754 156020
rect 508534 102704 511714 156020
rect 512494 102704 515434 156020
rect 516214 102704 519154 156020
rect 519934 102704 522874 156020
rect 523654 102704 526594 156020
rect 527374 102704 530314 156020
rect 482494 102580 530314 102704
rect 531094 102580 534034 156144
rect 534814 102580 537754 156144
rect 538534 102704 541714 156144
rect 542494 102704 552874 156144
rect 538534 102580 552874 102704
rect 553654 102580 556594 156144
rect 557374 102580 558676 156144
rect 456214 18144 558676 102580
rect 456214 8195 459154 18144
rect 459934 8195 462874 18144
rect 463654 8195 466594 18144
rect 467374 18020 485434 18144
rect 467374 8195 481714 18020
rect 482494 8195 485434 18020
rect 486214 18020 541714 18144
rect 486214 8195 489154 18020
rect 489934 8195 492874 18020
rect 493654 8195 496594 18020
rect 497374 8195 511714 18020
rect 512494 8195 515434 18020
rect 516214 8195 519154 18020
rect 519934 8195 522874 18020
rect 523654 8195 526594 18020
rect 527374 8195 541714 18020
rect 542494 18020 549154 18144
rect 542494 8195 545434 18020
rect 546214 8195 549154 18020
rect 549934 8195 552874 18144
rect 553654 8195 556594 18144
rect 557374 8195 558676 18144
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 700306 592650 700926
rect -8726 696586 592650 697206
rect -8726 692866 592650 693486
rect -8726 688906 592650 689526
rect -8726 685186 592650 685806
rect -8726 681466 592650 682086
rect -8726 677746 592650 678366
rect -8726 674026 592650 674646
rect -8726 670306 592650 670926
rect -8726 666586 592650 667206
rect -8726 662866 592650 663486
rect -8726 658906 592650 659526
rect -8726 655186 592650 655806
rect -8726 651466 592650 652086
rect -8726 647746 592650 648366
rect -8726 644026 592650 644646
rect -8726 640306 592650 640926
rect -8726 636586 592650 637206
rect -8726 632866 592650 633486
rect -8726 628906 592650 629526
rect -8726 625186 592650 625806
rect -8726 621466 592650 622086
rect -8726 617746 592650 618366
rect -8726 614026 592650 614646
rect -8726 610306 592650 610926
rect -8726 606586 592650 607206
rect -8726 602866 592650 603486
rect -8726 598906 592650 599526
rect -8726 595186 592650 595806
rect -8726 591466 592650 592086
rect -8726 587746 592650 588366
rect -8726 584026 592650 584646
rect -8726 580306 592650 580926
rect -8726 576586 592650 577206
rect -8726 572866 592650 573486
rect -8726 568906 592650 569526
rect -8726 565186 592650 565806
rect -8726 561466 592650 562086
rect -8726 557746 592650 558366
rect -8726 554026 592650 554646
rect -8726 550306 592650 550926
rect -8726 546586 592650 547206
rect -8726 542866 592650 543486
rect -8726 538906 592650 539526
rect -8726 535186 592650 535806
rect -8726 531466 592650 532086
rect -8726 527746 592650 528366
rect -8726 524026 592650 524646
rect -8726 520306 592650 520926
rect -8726 516586 592650 517206
rect -8726 512866 592650 513486
rect -8726 508906 592650 509526
rect -8726 505186 592650 505806
rect -8726 501466 592650 502086
rect -8726 497746 592650 498366
rect -8726 494026 592650 494646
rect -8726 490306 592650 490926
rect -8726 486586 592650 487206
rect -8726 482866 592650 483486
rect -8726 478906 592650 479526
rect -8726 475186 592650 475806
rect -8726 471466 592650 472086
rect -8726 467746 592650 468366
rect -8726 464026 592650 464646
rect -8726 460306 592650 460926
rect -8726 456586 592650 457206
rect -8726 452866 592650 453486
rect -8726 448906 592650 449526
rect -8726 445186 592650 445806
rect -8726 441466 592650 442086
rect -8726 437746 592650 438366
rect -8726 434026 592650 434646
rect -8726 430306 592650 430926
rect -8726 426586 592650 427206
rect -8726 422866 592650 423486
rect -8726 418906 592650 419526
rect -8726 415186 592650 415806
rect -8726 411466 592650 412086
rect -8726 407746 592650 408366
rect -8726 404026 592650 404646
rect -8726 400306 592650 400926
rect -8726 396586 592650 397206
rect -8726 392866 592650 393486
rect -8726 388906 592650 389526
rect -8726 385186 592650 385806
rect -8726 381466 592650 382086
rect -8726 377746 592650 378366
rect -8726 374026 592650 374646
rect -8726 370306 592650 370926
rect -8726 366586 592650 367206
rect -8726 362866 592650 363486
rect -8726 358906 592650 359526
rect -8726 355186 592650 355806
rect -8726 351466 592650 352086
rect -8726 347746 592650 348366
rect -8726 344026 592650 344646
rect -8726 340306 592650 340926
rect -8726 336586 592650 337206
rect -8726 332866 592650 333486
rect -8726 328906 592650 329526
rect -8726 325186 592650 325806
rect -8726 321466 592650 322086
rect -8726 317746 592650 318366
rect -8726 314026 592650 314646
rect -8726 310306 592650 310926
rect -8726 306586 592650 307206
rect -8726 302866 592650 303486
rect -8726 298906 592650 299526
rect -8726 295186 592650 295806
rect -8726 291466 592650 292086
rect -8726 287746 592650 288366
rect -8726 284026 592650 284646
rect -8726 280306 592650 280926
rect -8726 276586 592650 277206
rect -8726 272866 592650 273486
rect -8726 268906 592650 269526
rect -8726 265186 592650 265806
rect -8726 261466 592650 262086
rect -8726 257746 592650 258366
rect -8726 254026 592650 254646
rect -8726 250306 592650 250926
rect -8726 246586 592650 247206
rect -8726 242866 592650 243486
rect -8726 238906 592650 239526
rect -8726 235186 592650 235806
rect -8726 231466 592650 232086
rect -8726 227746 592650 228366
rect -8726 224026 592650 224646
rect -8726 220306 592650 220926
rect -8726 216586 592650 217206
rect -8726 212866 592650 213486
rect -8726 208906 592650 209526
rect -8726 205186 592650 205806
rect -8726 201466 592650 202086
rect -8726 197746 592650 198366
rect -8726 194026 592650 194646
rect -8726 190306 592650 190926
rect -8726 186586 592650 187206
rect -8726 182866 592650 183486
rect -8726 178906 592650 179526
rect -8726 175186 592650 175806
rect -8726 171466 592650 172086
rect -8726 167746 592650 168366
rect -8726 164026 592650 164646
rect -8726 160306 592650 160926
rect -8726 156586 592650 157206
rect -8726 152866 592650 153486
rect -8726 148906 592650 149526
rect -8726 145186 592650 145806
rect -8726 141466 592650 142086
rect -8726 137746 592650 138366
rect -8726 134026 592650 134646
rect -8726 130306 592650 130926
rect -8726 126586 592650 127206
rect -8726 122866 592650 123486
rect -8726 118906 592650 119526
rect -8726 115186 592650 115806
rect -8726 111466 592650 112086
rect -8726 107746 592650 108366
rect -8726 104026 592650 104646
rect -8726 100306 592650 100926
rect -8726 96586 592650 97206
rect -8726 92866 592650 93486
rect -8726 88906 592650 89526
rect -8726 85186 592650 85806
rect -8726 81466 592650 82086
rect -8726 77746 592650 78366
rect -8726 74026 592650 74646
rect -8726 70306 592650 70926
rect -8726 66586 592650 67206
rect -8726 62866 592650 63486
rect -8726 58906 592650 59526
rect -8726 55186 592650 55806
rect -8726 51466 592650 52086
rect -8726 47746 592650 48366
rect -8726 44026 592650 44646
rect -8726 40306 592650 40926
rect -8726 36586 592650 37206
rect -8726 32866 592650 33486
rect -8726 28906 592650 29526
rect -8726 25186 592650 25806
rect -8726 21466 592650 22086
rect -8726 17746 592650 18366
rect -8726 14026 592650 14646
rect -8726 10306 592650 10926
rect -8726 6586 592650 7206
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 31794 -7654 32414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 -7654 62414 17940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 102660 62414 155940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 240660 62414 293940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 378660 62414 423940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 508660 62414 569940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 61794 654660 62414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 -7654 92414 17940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 102784 92414 155940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 240784 92414 293940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 378784 92414 423940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 508784 92414 569940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 91794 654784 92414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 -7654 122414 18064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 102784 122414 156064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 240784 122414 294064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 378784 122414 424064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 508784 122414 570064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 121794 654784 122414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 151794 -7654 152414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 19199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 84857 182414 140559 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 654660 182414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 211794 -7654 212414 19199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 211794 84857 212414 140559 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 241794 -7654 242414 19199 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 241794 84857 242414 140559 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 241794 654784 242414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271794 -7654 272414 140559 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 271794 654784 272414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 301794 -7654 302414 140559 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 301794 539417 302414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 331794 -7654 332414 18064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 331794 654660 332414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 18064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 654784 362414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 391794 -7654 392414 18064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 391794 654660 392414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 421794 -7654 422414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 451794 -7654 452414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 -7654 482414 17940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 102660 482414 155940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 240660 482414 293940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 378660 482414 423940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 508660 482414 569940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 481794 654660 482414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 -7654 512414 17940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 102784 512414 155940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 240784 512414 293940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 378784 512414 423940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 508784 512414 569940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 511794 654784 512414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 18064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 102784 542414 156064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 240784 542414 294064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 378784 542414 424064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 508784 542414 570064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 654784 542414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 571794 -7654 572414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 32866 592650 33486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 62866 592650 63486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 92866 592650 93486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 122866 592650 123486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 152866 592650 153486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 212866 592650 213486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 242866 592650 243486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 272866 592650 273486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 302866 592650 303486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 332866 592650 333486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 392866 592650 393486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 422866 592650 423486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 452866 592650 453486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 482866 592650 483486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 512866 592650 513486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 572866 592650 573486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 602866 592650 603486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 632866 592650 633486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 662866 592650 663486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 692866 592650 693486 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 9234 -7654 9854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 39234 -7654 39854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 39234 240660 39854 294064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 39234 508660 39854 570064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 39234 654660 39854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 -7654 69854 17940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 102784 69854 155940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 240784 69854 293940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 378784 69854 423940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 508784 69854 569940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 69234 654784 69854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 -7654 99854 17940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 102784 99854 155940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 240784 99854 293940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 378784 99854 423940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 508784 99854 569940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 99234 654784 99854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 129234 -7654 129854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 129234 240660 129854 294064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 129234 508660 129854 570064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 129234 654660 129854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 159234 -7654 159854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 -7654 189854 19199 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 84857 189854 140559 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 654660 189854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219234 -7654 219854 19199 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219234 84857 219854 140559 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219234 654784 219854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 249234 -7654 249854 19199 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 249234 84857 249854 140559 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 249234 654660 249854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 279234 -7654 279854 140559 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 279234 654660 279854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 309234 -7654 309854 140559 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 309234 539417 309854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 339234 -7654 339854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 339234 654660 339854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 -7654 369854 17940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 654784 369854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 399234 -7654 399854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 399234 654660 399854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 429234 -7654 429854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 459234 -7654 459854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 459234 240660 459854 294064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 459234 508660 459854 570064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 459234 654660 459854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 -7654 489854 17940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 102784 489854 155940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 240784 489854 293940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 378784 489854 423940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 508784 489854 569940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 489234 654784 489854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 -7654 519854 17940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 102784 519854 155940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 240784 519854 293940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 378784 519854 423940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 508784 519854 569940 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 519234 654784 519854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 -7654 549854 18064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 240660 549854 294064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 508660 549854 570064 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 654660 549854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 579234 -7654 579854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 10306 592650 10926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 40306 592650 40926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 70306 592650 70926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 100306 592650 100926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 130306 592650 130926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 160306 592650 160926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 190306 592650 190926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 220306 592650 220926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 250306 592650 250926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 280306 592650 280926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 310306 592650 310926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 340306 592650 340926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 370306 592650 370926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 400306 592650 400926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 430306 592650 430926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 460306 592650 460926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 490306 592650 490926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 520306 592650 520926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 550306 592650 550926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 580306 592650 580926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 610306 592650 610926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 640306 592650 640926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 670306 592650 670926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 700306 592650 700926 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 16674 -7654 17294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46674 -7654 47294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46674 102660 47294 156064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46674 240660 47294 294064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46674 508660 47294 570064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 46674 654660 47294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 -7654 77294 17940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 102784 77294 155940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 240784 77294 293940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 378784 77294 423940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 508784 77294 569940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 76674 654784 77294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 -7654 107294 17940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 102784 107294 155940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 240784 107294 293940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 378784 107294 423940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 508784 107294 569940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 106674 654784 107294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136674 -7654 137294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136674 102660 137294 156064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136674 240660 137294 294064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136674 508660 137294 570064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 136674 654660 137294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 166674 -7654 167294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 -7654 197294 19199 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 84857 197294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 654660 197294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 226674 -7654 227294 19199 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 226674 84857 227294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 256674 -7654 257294 19199 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 256674 84857 257294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 256674 654660 257294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 286674 -7654 287294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 286674 539417 287294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 316674 -7654 317294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 316674 539417 317294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 346674 -7654 347294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 346674 102660 347294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 346674 654660 347294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 -7654 377294 17940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 102784 377294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 654784 377294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 406674 -7654 407294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 406674 102660 407294 140559 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 406674 654660 407294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 436674 -7654 437294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 466674 -7654 467294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 466674 102660 467294 156064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 466674 240660 467294 294064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 466674 508660 467294 570064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 466674 654660 467294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 -7654 497294 17940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 102784 497294 155940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 240784 497294 293940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 378784 497294 423940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 508784 497294 569940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 496674 654784 497294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 -7654 527294 17940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 102784 527294 155940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 240784 527294 293940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 378784 527294 423940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 508784 527294 569940 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 526674 654784 527294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 -7654 557294 18064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 102660 557294 156064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 240660 557294 294064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 508660 557294 570064 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 654660 557294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 17746 592650 18366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 47746 592650 48366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 77746 592650 78366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 107746 592650 108366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 137746 592650 138366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 167746 592650 168366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 197746 592650 198366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 227746 592650 228366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 257746 592650 258366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 287746 592650 288366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 317746 592650 318366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 347746 592650 348366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 377746 592650 378366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 407746 592650 408366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 437746 592650 438366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 467746 592650 468366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 497746 592650 498366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 527746 592650 528366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 557746 592650 558366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 587746 592650 588366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 617746 592650 618366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 647746 592650 648366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 677746 592650 678366 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 24114 -7654 24734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54114 102660 54734 156064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54114 378660 54734 424064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54114 508660 54734 570064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 54114 654660 54734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84114 102784 84734 155940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84114 240784 84734 293940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84114 378784 84734 423940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84114 508784 84734 569940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 84114 654784 84734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 114114 102660 114734 156064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 114114 378660 114734 424064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 114114 508660 114734 570064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 114114 654660 114734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 144114 -7654 144734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 174114 -7654 174734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 84857 204734 140559 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 654660 204734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 234114 84857 234734 140559 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 234114 654784 234734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 264114 84857 264734 140559 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 264114 654660 264734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 294114 -7654 294734 140559 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 294114 539417 294734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 324114 654660 324734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 354114 654784 354734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 654784 384734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 414114 654660 414734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 444114 -7654 444734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474114 102660 474734 156064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474114 378660 474734 424064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474114 508660 474734 570064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 474114 654660 474734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 504114 102784 504734 155940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 504114 240784 504734 293940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 504114 378784 504734 423940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 504114 508784 504734 569940 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 504114 654784 504734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 534114 102660 534734 156064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 534114 378660 534734 424064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 534114 508660 534734 570064 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 534114 654660 534734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 564114 -7654 564734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 25186 592650 25806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 55186 592650 55806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 85186 592650 85806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 115186 592650 115806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 145186 592650 145806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 175186 592650 175806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 205186 592650 205806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 235186 592650 235806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 265186 592650 265806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 295186 592650 295806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 325186 592650 325806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 355186 592650 355806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 385186 592650 385806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 415186 592650 415806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 445186 592650 445806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 475186 592650 475806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 505186 592650 505806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 535186 592650 535806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 565186 592650 565806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 595186 592650 595806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 625186 592650 625806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 655186 592650 655806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 685186 592650 685806 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 20394 -7654 21014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 50394 102660 51014 156064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 50394 240660 51014 294064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 50394 378660 51014 424064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 50394 508660 51014 570064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 50394 654660 51014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 80394 102784 81014 155940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 80394 240784 81014 293940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 80394 378784 81014 423940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 80394 508784 81014 569940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 80394 654784 81014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 110394 102660 111014 156064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 110394 240660 111014 294064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 110394 378660 111014 424064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 110394 508660 111014 570064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 110394 654660 111014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 140394 -7654 141014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 170394 -7654 171014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 654660 201014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 230394 654784 231014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 260394 654660 261014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 290394 -7654 291014 140559 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 290394 539417 291014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 320394 654784 321014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 350394 654784 351014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 654784 381014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 410394 654660 411014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 440394 -7654 441014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 470394 102660 471014 156064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 470394 240660 471014 294064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 470394 378660 471014 424064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 470394 508660 471014 570064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 470394 654660 471014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 500394 102784 501014 155940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 500394 240784 501014 293940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 500394 378784 501014 423940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 500394 508784 501014 569940 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 500394 654784 501014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 530394 102660 531014 156064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 530394 240660 531014 294064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 530394 378660 531014 424064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 530394 508660 531014 570064 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 530394 654660 531014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 560394 -7654 561014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 21466 592650 22086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 51466 592650 52086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 81466 592650 82086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 111466 592650 112086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 141466 592650 142086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 171466 592650 172086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 201466 592650 202086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 231466 592650 232086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 261466 592650 262086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 291466 592650 292086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 321466 592650 322086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 351466 592650 352086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 381466 592650 382086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 411466 592650 412086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 441466 592650 442086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 471466 592650 472086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 501466 592650 502086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 531466 592650 532086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 561466 592650 562086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 591466 592650 592086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 621466 592650 622086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 651466 592650 652086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 681466 592650 682086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 27834 -7654 28454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 57834 102660 58454 155940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 57834 378660 58454 423940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 57834 508660 58454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 57834 654660 58454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 87834 102784 88454 155940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 87834 240784 88454 293940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 87834 378784 88454 423940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 87834 508784 88454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 87834 654784 88454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 117834 102660 118454 156064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 117834 378660 118454 424064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 117834 508660 118454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 117834 654660 118454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 147834 -7654 148454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 177834 -7654 178454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 177834 654660 178454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 84857 208454 140559 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 539417 208454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 654660 208454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 237834 84857 238454 140559 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 237834 539417 238454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 237834 654784 238454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 267834 84857 268454 140559 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 267834 539417 268454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 267834 654660 268454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 297834 -7654 298454 140559 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 297834 539417 298454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 327834 539417 328454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 327834 654660 328454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 357834 539417 358454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 357834 654784 358454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 539417 388454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 654784 388454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 417834 539417 418454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 417834 654784 418454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 447834 -7654 448454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477834 102660 478454 155940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477834 378660 478454 423940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477834 508660 478454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477834 654660 478454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 507834 102784 508454 155940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 507834 240784 508454 293940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 507834 378784 508454 423940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 507834 508784 508454 569940 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 507834 654784 508454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 537834 102660 538454 156064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 537834 378660 538454 424064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 537834 508660 538454 570064 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 537834 654660 538454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 567834 -7654 568454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 28906 592650 29526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 58906 592650 59526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 88906 592650 89526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 118906 592650 119526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 148906 592650 149526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 178906 592650 179526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 208906 592650 209526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 238906 592650 239526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 268906 592650 269526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 298906 592650 299526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 328906 592650 329526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 358906 592650 359526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 388906 592650 389526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 418906 592650 419526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 448906 592650 449526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 478906 592650 479526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 508906 592650 509526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 538906 592650 539526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 568906 592650 569526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 598906 592650 599526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 628906 592650 629526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 658906 592650 659526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 688906 592650 689526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 5514 -7654 6134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 35514 -7654 36134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65514 -7654 66134 18064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65514 240660 66134 294064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65514 508660 66134 570064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65514 654660 66134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 -7654 96134 17940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 102784 96134 155940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 240784 96134 293940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 378784 96134 423940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 508784 96134 569940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 95514 654784 96134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 125514 -7654 126134 17940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 125514 240660 126134 293940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 125514 508660 126134 569940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 125514 654660 126134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 155514 -7654 156134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 -7654 186134 19199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 84857 186134 140559 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 654660 186134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 215514 -7654 216134 19199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 215514 84857 216134 140559 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 215514 654784 216134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 245514 -7654 246134 19199 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 245514 654784 246134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 275514 -7654 276134 140559 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 275514 654660 276134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 305514 -7654 306134 140559 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 305514 539417 306134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 335514 -7654 336134 18064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 335514 654660 336134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 -7654 366134 17940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 654784 366134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 395514 -7654 396134 18064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 395514 654660 396134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 425514 -7654 426134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 455514 -7654 456134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485514 -7654 486134 18064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485514 240660 486134 294064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485514 508660 486134 570064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 485514 654660 486134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 -7654 516134 17940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 102784 516134 155940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 240784 516134 293940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 378784 516134 423940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 508784 516134 569940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 515514 654784 516134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 -7654 546134 17940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 240660 546134 293940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 508660 546134 569940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 654660 546134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 575514 -7654 576134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 6586 592650 7206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 36586 592650 37206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 66586 592650 67206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 96586 592650 97206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 126586 592650 127206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 156586 592650 157206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 186586 592650 187206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 216586 592650 217206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 246586 592650 247206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 276586 592650 277206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 306586 592650 307206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 336586 592650 337206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 366586 592650 367206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 396586 592650 397206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 426586 592650 427206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 456586 592650 457206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 486586 592650 487206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 516586 592650 517206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 546586 592650 547206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 576586 592650 577206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 606586 592650 607206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 636586 592650 637206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 666586 592650 667206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 696586 592650 697206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42954 -7654 43574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42954 102660 43574 156064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42954 240660 43574 294064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42954 508660 43574 570064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 42954 654660 43574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 -7654 73574 17940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 102784 73574 155940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 240784 73574 293940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 378784 73574 423940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 508784 73574 569940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 72954 654784 73574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 -7654 103574 17940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 102784 103574 155940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 240784 103574 293940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 378784 103574 423940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 508784 103574 569940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 102954 654784 103574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132954 -7654 133574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132954 102660 133574 156064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132954 240660 133574 294064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132954 508660 133574 570064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 132954 654660 133574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 162954 -7654 163574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 -7654 193574 19199 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 84857 193574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 654660 193574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222954 -7654 223574 19199 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222954 84857 223574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222954 654784 223574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 252954 -7654 253574 19199 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 252954 84857 253574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 252954 654660 253574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 282954 -7654 283574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 282954 539417 283574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 312954 -7654 313574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 312954 539417 313574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 342954 -7654 343574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 342954 102660 343574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 342954 654660 343574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 -7654 373574 17940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 102784 373574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 654784 373574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 402954 -7654 403574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 402954 102784 403574 140559 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 402954 654660 403574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 432954 -7654 433574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 462954 -7654 463574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 462954 102660 463574 156064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 462954 240660 463574 294064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 462954 508660 463574 570064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 462954 654660 463574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 -7654 493574 17940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 102784 493574 155940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 240784 493574 293940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 378784 493574 423940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 508784 493574 569940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 492954 654784 493574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 -7654 523574 17940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 102784 523574 155940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 240784 523574 293940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 378784 523574 423940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 508784 523574 569940 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 522954 654784 523574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 -7654 553574 18064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 102660 553574 156064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 240660 553574 294064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 508660 553574 570064 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 654660 553574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 44026 592650 44646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 74026 592650 74646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 104026 592650 104646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 134026 592650 134646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 164026 592650 164646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 224026 592650 224646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 254026 592650 254646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 284026 592650 284646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 314026 592650 314646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 344026 592650 344646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 404026 592650 404646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 434026 592650 434646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 464026 592650 464646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 494026 592650 494646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 524026 592650 524646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 584026 592650 584646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 614026 592650 614646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 644026 592650 644646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 674026 592650 674646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 291914412
string GDS_FILE /home/tobi/proj/STW/8c/stw_8c_release/STW_8/openlane/user_project_wrapper/runs/22_12_10_07_53/results/signoff/user_project_wrapper.magic.gds
string GDS_START 286244558
<< end >>

